
module fp_1 ( clock, reset, in1, in2, in3, in4, ops_out );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  output [31:0] ops_out;
  input clock, reset;
  wire   U6_Z_0, U6_Z_1, U6_Z_2, U6_Z_3, U6_Z_4, U6_Z_5, U6_Z_6, U6_Z_7,
         U6_Z_8, U6_Z_9, U6_Z_10, U6_Z_11, U6_Z_12, U6_Z_13, U6_Z_14, U6_Z_15,
         U6_Z_16, U6_Z_17, U6_Z_18, U6_Z_19, U6_Z_20, U6_Z_21, U6_Z_22,
         U6_Z_23, U6_Z_24, U6_Z_25, U6_Z_26, U6_Z_27, U6_Z_28, U6_Z_29,
         U6_Z_30, U6_Z_31, U5_Z_0, U5_Z_1, U5_Z_2, U5_Z_3, U5_Z_4, U5_Z_5,
         U5_Z_6, U5_Z_7, U5_Z_8, U5_Z_9, U5_Z_10, U5_Z_11, U5_Z_12, U5_Z_13,
         U5_Z_14, U5_Z_15, U5_Z_16, U5_Z_17, U5_Z_18, U5_Z_19, U5_Z_20,
         U5_Z_21, U5_Z_22, U5_Z_23, U5_Z_24, U5_Z_25, U5_Z_26, U5_Z_27,
         U5_Z_28, U5_Z_29, U5_Z_30, U5_Z_31, U4_Z_1, U4_Z_2, U4_Z_3, U4_Z_4,
         U4_Z_5, U4_Z_6, U4_Z_7, U4_Z_8, U4_Z_9, U4_Z_10, U4_Z_11, U4_Z_12,
         U4_Z_13, U4_Z_14, U4_Z_15, U4_Z_16, U4_Z_17, U4_Z_18, U4_Z_19,
         U4_Z_20, U4_Z_21, U4_Z_22, U4_Z_23, U4_Z_24, U4_Z_25, U4_Z_26,
         U4_Z_27, U4_Z_28, U4_Z_29, U4_Z_30, U4_Z_31, add_49_B_0_, add_49_B_1_,
         add_49_B_2_, add_49_B_3_, add_49_B_4_, add_49_B_5_, add_49_B_6_,
         add_49_B_7_, add_49_B_8_, add_49_B_9_, add_49_B_10_, add_49_B_11_,
         add_49_B_12_, add_49_B_13_, add_49_B_14_, add_49_B_15_, add_49_B_16_,
         add_49_B_17_, add_49_B_18_, add_49_B_19_, add_49_B_20_, add_49_B_21_,
         add_49_B_22_, add_49_B_23_, add_49_B_24_, add_49_B_25_, add_49_B_26_,
         add_49_B_27_, add_49_B_28_, add_49_B_29_, add_49_B_30_, add_49_B_31_,
         add_49_A_0_, add_49_A_1_, add_49_A_2_, add_49_A_3_, add_49_A_4_,
         add_49_A_5_, add_49_A_6_, add_49_A_7_, add_49_A_8_, add_49_A_9_,
         add_49_A_10_, add_49_A_11_, add_49_A_12_, add_49_A_13_, add_49_A_14_,
         add_49_A_15_, add_49_A_16_, add_49_A_17_, add_49_A_18_, add_49_A_19_,
         add_49_A_20_, add_49_A_21_, add_49_A_22_, add_49_A_23_, add_49_A_24_,
         add_49_A_25_, add_49_A_26_, add_49_A_27_, add_49_A_28_, add_49_A_29_,
         add_49_A_30_, add_49_A_31_, net1690, net1701, net1703, net1722,
         net1724, net1726, net1727, net1750, net1751, net1798, net1815,
         net1817, net1818, net1855, net1861, net2053, net2094, net2119,
         net2123, net2125, net2175, net2177, net2188, net2213, net2222,
         net2399, net2489, net2482, net2513, net2722, net2804, net2805,
         net2879, net2882, net2902, net2982, net3004, net3065, net3098,
         net3132, net3189, net3196, net3406, net3421, net3443, net3442,
         net3455, net3472, net3479, net3503, net3542, net3768, net3757,
         net3979, net3978, net4289, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226;

  DFF_X2 adr_2_op_reg_30_ ( .D(U4_Z_30), .CK(clock), .Q(add_49_B_30_), .QN(
        n1222) );
  DFF_X2 adr_2_op_reg_0_ ( .D(n862), .CK(clock), .Q(add_49_B_0_) );
  DFF_X2 adr_1_op_reg_0_ ( .D(U5_Z_0), .CK(clock), .Q(add_49_A_0_) );
  DFF_X2 adr_1_op_reg_1_ ( .D(U5_Z_1), .CK(clock), .Q(add_49_A_1_), .QN(n904)
         );
  DFF_X2 adr_2_op_reg_3_ ( .D(U4_Z_3), .CK(clock), .Q(add_49_B_3_), .QN(n538)
         );
  DFF_X2 adr_2_op_reg_2_ ( .D(U4_Z_2), .CK(clock), .Q(add_49_B_2_), .QN(n920)
         );
  DFF_X2 adr_2_op_reg_1_ ( .D(U4_Z_1), .CK(clock), .Q(add_49_B_1_), .QN(n903)
         );
  DFF_X2 adr_1_op_reg_2_ ( .D(U5_Z_2), .CK(clock), .Q(add_49_A_2_), .QN(n921)
         );
  DFF_X2 adr_2_op_reg_4_ ( .D(U4_Z_4), .CK(clock), .Q(add_49_B_4_), .QN(n953)
         );
  DFF_X2 adr_1_op_reg_3_ ( .D(U5_Z_3), .CK(clock), .Q(add_49_A_3_), .QN(n539)
         );
  DFF_X2 adr_2_op_reg_5_ ( .D(U4_Z_5), .CK(clock), .Q(add_49_B_5_) );
  DFF_X2 adr_1_op_reg_4_ ( .D(U5_Z_4), .CK(clock), .Q(add_49_A_4_), .QN(n954)
         );
  DFF_X2 adr_1_op_reg_5_ ( .D(U5_Z_5), .CK(clock), .Q(add_49_A_5_) );
  DFF_X2 adr_2_op_reg_7_ ( .D(U4_Z_7), .CK(clock), .Q(add_49_B_7_), .QN(n996)
         );
  DFF_X2 adr_2_op_reg_6_ ( .D(U4_Z_6), .CK(clock), .Q(add_49_B_6_), .QN(n982)
         );
  DFF_X2 adr_2_op_reg_8_ ( .D(U4_Z_8), .CK(clock), .Q(add_49_B_8_), .QN(n1011)
         );
  DFF_X2 adr_1_op_reg_6_ ( .D(U5_Z_6), .CK(clock), .Q(add_49_A_6_), .QN(n983)
         );
  DFF_X2 adr_2_op_reg_9_ ( .D(U4_Z_9), .CK(clock), .Q(add_49_B_9_), .QN(n536)
         );
  DFF_X2 adr_1_op_reg_7_ ( .D(U5_Z_7), .CK(clock), .Q(add_49_A_7_), .QN(n997)
         );
  DFF_X2 adr_1_op_reg_8_ ( .D(U5_Z_8), .CK(clock), .Q(add_49_A_8_), .QN(n1012)
         );
  DFF_X2 adr_2_op_reg_10_ ( .D(U4_Z_10), .CK(clock), .Q(add_49_B_10_), .QN(
        n1034) );
  DFF_X2 adr_2_op_reg_11_ ( .D(U4_Z_11), .CK(clock), .Q(add_49_B_11_), .QN(
        n546) );
  DFF_X2 adr_1_op_reg_10_ ( .D(U5_Z_10), .CK(clock), .Q(add_49_A_10_), .QN(
        n1035) );
  DFF_X2 adr_1_op_reg_9_ ( .D(U5_Z_9), .CK(clock), .Q(add_49_A_9_), .QN(n537)
         );
  DFF_X2 adr_2_op_reg_12_ ( .D(U4_Z_12), .CK(clock), .Q(add_49_B_12_), .QN(
        n1053) );
  DFF_X2 adr_1_op_reg_11_ ( .D(U5_Z_11), .CK(clock), .Q(add_49_A_11_), .QN(
        n547) );
  DFF_X2 adr_1_op_reg_12_ ( .D(U5_Z_12), .CK(clock), .Q(add_49_A_12_), .QN(
        n1054) );
  DFF_X2 adr_1_op_reg_13_ ( .D(U5_Z_13), .CK(clock), .Q(add_49_A_13_), .QN(
        n530) );
  DFF_X2 adr_2_op_reg_13_ ( .D(U4_Z_13), .CK(clock), .Q(add_49_B_13_), .QN(
        n529) );
  DFF_X2 adr_2_op_reg_14_ ( .D(U4_Z_14), .CK(clock), .Q(add_49_B_14_), .QN(
        n1069) );
  DFF_X2 adr_1_op_reg_14_ ( .D(U5_Z_14), .CK(clock), .Q(add_49_A_14_), .QN(
        n1070) );
  DFF_X2 adr_1_op_reg_15_ ( .D(U5_Z_15), .CK(clock), .Q(add_49_A_15_), .QN(
        n535) );
  DFF_X2 adr_1_op_reg_16_ ( .D(U5_Z_16), .CK(clock), .Q(add_49_A_16_), .QN(
        n1089) );
  DFF_X2 adr_2_op_reg_15_ ( .D(U4_Z_15), .CK(clock), .Q(add_49_B_15_), .QN(
        n534) );
  DFF_X2 adr_1_op_reg_17_ ( .D(U5_Z_17), .CK(clock), .Q(add_49_A_17_), .QN(
        n551) );
  DFF_X2 adr_2_op_reg_16_ ( .D(U4_Z_16), .CK(clock), .Q(add_49_B_16_), .QN(
        n1088) );
  DFF_X2 adr_1_op_reg_18_ ( .D(U5_Z_18), .CK(clock), .Q(add_49_A_18_), .QN(
        n1111) );
  DFF_X2 adr_2_op_reg_17_ ( .D(U4_Z_17), .CK(clock), .Q(add_49_B_17_), .QN(
        n550) );
  DFF_X2 adr_1_op_reg_19_ ( .D(U5_Z_19), .CK(clock), .Q(add_49_A_19_), .QN(
        n545) );
  DFF_X2 adr_2_op_reg_18_ ( .D(U4_Z_18), .CK(clock), .Q(add_49_B_18_), .QN(
        n1110) );
  DFF_X2 adr_1_op_reg_20_ ( .D(U5_Z_20), .CK(clock), .Q(add_49_A_20_), .QN(
        n1142) );
  DFF_X2 adr_2_op_reg_19_ ( .D(U4_Z_19), .CK(clock), .Q(add_49_B_19_), .QN(
        n544) );
  DFF_X2 adr_2_op_reg_20_ ( .D(U4_Z_20), .CK(clock), .Q(add_49_B_20_), .QN(
        n1141) );
  DFF_X2 adr_1_op_reg_21_ ( .D(U5_Z_21), .CK(clock), .Q(add_49_A_21_), .QN(
        n533) );
  DFF_X2 adr_2_op_reg_21_ ( .D(U4_Z_21), .CK(clock), .Q(add_49_B_21_), .QN(
        n532) );
  DFF_X2 adr_1_op_reg_22_ ( .D(U5_Z_22), .CK(clock), .Q(add_49_A_22_), .QN(
        n1168) );
  DFF_X2 adr_1_op_reg_23_ ( .D(U5_Z_23), .CK(clock), .Q(add_49_A_23_), .QN(
        n528) );
  DFF_X2 adr_2_op_reg_22_ ( .D(U4_Z_22), .CK(clock), .Q(add_49_B_22_), .QN(
        n1167) );
  DFF_X2 adr_1_op_reg_24_ ( .D(U5_Z_24), .CK(clock), .Q(add_49_A_24_), .QN(
        n1185) );
  DFF_X2 adr_2_op_reg_23_ ( .D(U4_Z_23), .CK(clock), .Q(add_49_B_23_), .QN(
        n527) );
  DFF_X2 adr_1_op_reg_25_ ( .D(U5_Z_25), .CK(clock), .Q(add_49_A_25_), .QN(
        n543) );
  DFF_X2 adr_2_op_reg_24_ ( .D(U4_Z_24), .CK(clock), .Q(add_49_B_24_), .QN(
        n1184) );
  DFF_X2 adr_1_op_reg_27_ ( .D(U5_Z_27), .CK(clock), .Q(add_49_A_27_) );
  DFF_X2 adr_1_op_reg_26_ ( .D(U5_Z_26), .CK(clock), .Q(add_49_A_26_), .QN(
        n1202) );
  DFF_X2 adr_1_op_reg_28_ ( .D(U5_Z_28), .CK(clock), .Q(add_49_A_28_), .QN(
        n1214) );
  DFF_X2 adr_2_op_reg_27_ ( .D(U4_Z_27), .CK(clock), .Q(add_49_B_27_) );
  DFF_X2 adr_1_op_reg_29_ ( .D(U5_Z_29), .CK(clock), .Q(add_49_A_29_), .QN(
        n526) );
  DFF_X2 adr_1_op_reg_30_ ( .D(U5_Z_30), .CK(clock), .Q(add_49_A_30_), .QN(
        n1223) );
  DFF_X2 adr_2_op_reg_28_ ( .D(U4_Z_28), .CK(clock), .Q(add_49_B_28_), .QN(
        n1213) );
  DFF_X2 adr_2_op_reg_29_ ( .D(U4_Z_29), .CK(clock), .Q(add_49_B_29_), .QN(
        n525) );
  DFF_X2 ops_out_reg_0_ ( .D(U6_Z_0), .CK(clock), .Q(ops_out[0]) );
  DFF_X2 ops_out_reg_2_ ( .D(U6_Z_2), .CK(clock), .Q(ops_out[2]) );
  DFF_X2 ops_out_reg_1_ ( .D(U6_Z_1), .CK(clock), .Q(ops_out[1]) );
  DFF_X2 ops_out_reg_3_ ( .D(U6_Z_3), .CK(clock), .Q(ops_out[3]) );
  DFF_X2 ops_out_reg_4_ ( .D(U6_Z_4), .CK(clock), .Q(ops_out[4]) );
  DFF_X2 ops_out_reg_5_ ( .D(U6_Z_5), .CK(clock), .Q(ops_out[5]) );
  DFF_X2 ops_out_reg_6_ ( .D(U6_Z_6), .CK(clock), .Q(ops_out[6]) );
  DFF_X2 ops_out_reg_7_ ( .D(U6_Z_7), .CK(clock), .Q(ops_out[7]) );
  DFF_X2 ops_out_reg_8_ ( .D(U6_Z_8), .CK(clock), .Q(ops_out[8]) );
  DFF_X2 ops_out_reg_9_ ( .D(U6_Z_9), .CK(clock), .Q(ops_out[9]) );
  DFF_X2 ops_out_reg_10_ ( .D(U6_Z_10), .CK(clock), .Q(ops_out[10]) );
  DFF_X2 ops_out_reg_11_ ( .D(U6_Z_11), .CK(clock), .Q(ops_out[11]) );
  DFF_X2 ops_out_reg_12_ ( .D(U6_Z_12), .CK(clock), .Q(ops_out[12]) );
  DFF_X2 ops_out_reg_13_ ( .D(U6_Z_13), .CK(clock), .Q(ops_out[13]) );
  DFF_X2 ops_out_reg_14_ ( .D(U6_Z_14), .CK(clock), .Q(ops_out[14]) );
  DFF_X2 ops_out_reg_15_ ( .D(U6_Z_15), .CK(clock), .Q(ops_out[15]) );
  DFF_X2 ops_out_reg_16_ ( .D(U6_Z_16), .CK(clock), .Q(ops_out[16]) );
  DFF_X2 ops_out_reg_17_ ( .D(U6_Z_17), .CK(clock), .Q(ops_out[17]) );
  DFF_X2 ops_out_reg_18_ ( .D(U6_Z_18), .CK(clock), .Q(ops_out[18]) );
  DFF_X2 ops_out_reg_19_ ( .D(U6_Z_19), .CK(clock), .Q(ops_out[19]) );
  DFF_X2 ops_out_reg_20_ ( .D(U6_Z_20), .CK(clock), .Q(ops_out[20]) );
  DFF_X2 ops_out_reg_21_ ( .D(U6_Z_21), .CK(clock), .Q(ops_out[21]) );
  DFF_X2 ops_out_reg_22_ ( .D(U6_Z_22), .CK(clock), .Q(ops_out[22]) );
  DFF_X2 ops_out_reg_23_ ( .D(U6_Z_23), .CK(clock), .Q(ops_out[23]) );
  DFF_X2 ops_out_reg_24_ ( .D(U6_Z_24), .CK(clock), .Q(ops_out[24]) );
  DFF_X2 ops_out_reg_25_ ( .D(U6_Z_25), .CK(clock), .Q(ops_out[25]) );
  DFF_X2 ops_out_reg_26_ ( .D(U6_Z_26), .CK(clock), .Q(ops_out[26]) );
  DFF_X2 ops_out_reg_27_ ( .D(U6_Z_27), .CK(clock), .Q(ops_out[27]) );
  DFF_X2 ops_out_reg_28_ ( .D(U6_Z_28), .CK(clock), .Q(ops_out[28]) );
  DFF_X2 ops_out_reg_29_ ( .D(U6_Z_29), .CK(clock), .Q(ops_out[29]) );
  DFF_X2 ops_out_reg_30_ ( .D(U6_Z_30), .CK(clock), .Q(ops_out[30]) );
  DFF_X2 adr_2_op_reg_25_ ( .D(U4_Z_25), .CK(clock), .Q(add_49_B_25_), .QN(
        n542) );
  DFF_X2 adr_2_op_reg_26_ ( .D(U4_Z_26), .CK(clock), .Q(add_49_B_26_), .QN(
        n1201) );
  DFF_X2 adr_1_op_reg_31_ ( .D(U5_Z_31), .CK(clock), .Q(add_49_A_31_) );
  DFF_X2 ops_out_reg_31_ ( .D(U6_Z_31), .CK(clock), .Q(ops_out[31]) );
  DFF_X2 adr_2_op_reg_31_ ( .D(U4_Z_31), .CK(clock), .Q(add_49_B_31_) );
  NOR2_X4 U170 ( .A1(net2882), .A2(n660), .ZN(n596) );
  INV_X2 U171 ( .A(n779), .ZN(n549) );
  INV_X4 U172 ( .A(n747), .ZN(n1028) );
  NOR2_X4 U173 ( .A1(n747), .A2(n1030), .ZN(n741) );
  INV_X2 U174 ( .A(n548), .ZN(n678) );
  INV_X2 U175 ( .A(n686), .ZN(n687) );
  NOR2_X2 U176 ( .A1(n1161), .A2(n1162), .ZN(net3132) );
  NOR2_X2 U177 ( .A1(n732), .A2(n1084), .ZN(n743) );
  OR2_X4 U178 ( .A1(in2[0]), .A2(in4[29]), .ZN(n659) );
  AND2_X4 U179 ( .A1(n642), .A2(n618), .ZN(n531) );
  NAND2_X2 U180 ( .A1(n525), .A2(n526), .ZN(n591) );
  NAND2_X2 U181 ( .A1(n527), .A2(n528), .ZN(n581) );
  NAND2_X2 U182 ( .A1(n529), .A2(n530), .ZN(n571) );
  NAND2_X2 U183 ( .A1(n945), .A2(in4[4]), .ZN(n946) );
  OAI21_X2 U184 ( .B1(n792), .B2(in2[4]), .A(n713), .ZN(n898) );
  XNOR2_X1 U185 ( .A(n886), .B(in4[0]), .ZN(n881) );
  AND3_X4 U186 ( .A1(net1724), .A2(n654), .A3(n560), .ZN(n670) );
  NOR2_X2 U187 ( .A1(n1082), .A2(n1083), .ZN(n744) );
  OAI22_X2 U188 ( .A1(n806), .A2(n785), .B1(n1092), .B2(n784), .ZN(n567) );
  OAI22_X2 U189 ( .A1(n618), .A2(net1855), .B1(n531), .B2(n629), .ZN(net1818)
         );
  NAND2_X2 U190 ( .A1(n532), .A2(n533), .ZN(n577) );
  NAND2_X2 U191 ( .A1(n534), .A2(n535), .ZN(n572) );
  NAND2_X2 U192 ( .A1(n536), .A2(n537), .ZN(n570) );
  NAND2_X2 U193 ( .A1(n538), .A2(n539), .ZN(n564) );
  OAI22_X2 U194 ( .A1(in4[25]), .A2(in2[28]), .B1(in4[26]), .B2(in2[29]), .ZN(
        n627) );
  OAI21_X2 U195 ( .B1(n540), .B2(in3[12]), .A(n610), .ZN(n599) );
  INV_X4 U196 ( .A(net3768), .ZN(n540) );
  NAND3_X2 U197 ( .A1(n541), .A2(n668), .A3(n964), .ZN(n798) );
  INV_X4 U198 ( .A(in4[6]), .ZN(n541) );
  XNOR2_X2 U199 ( .A(in4[4]), .B(n948), .ZN(n935) );
  XNOR2_X2 U200 ( .A(in4[2]), .B(n916), .ZN(n899) );
  NAND3_X1 U201 ( .A1(n640), .A2(n636), .A3(net3421), .ZN(n644) );
  XNOR2_X2 U202 ( .A(in1[20]), .B(in1[18]), .ZN(n883) );
  NAND2_X2 U203 ( .A1(n542), .A2(n543), .ZN(n582) );
  NAND2_X2 U204 ( .A1(n544), .A2(n545), .ZN(n576) );
  NAND2_X2 U205 ( .A1(n546), .A2(n547), .ZN(n569) );
  AOI21_X2 U206 ( .B1(n618), .B2(n642), .A(n629), .ZN(n625) );
  OAI21_X1 U207 ( .B1(n597), .B2(n1059), .A(n719), .ZN(n548) );
  NAND3_X2 U208 ( .A1(net3768), .A2(n693), .A3(n692), .ZN(n698) );
  OAI22_X2 U209 ( .A1(n674), .A2(n1006), .B1(n1008), .B2(n1007), .ZN(n675) );
  XNOR2_X2 U210 ( .A(n949), .B(in2[8]), .ZN(n563) );
  NAND3_X1 U211 ( .A1(n791), .A2(n790), .A3(in2[3]), .ZN(n787) );
  XNOR2_X1 U212 ( .A(n930), .B(n917), .ZN(n918) );
  NOR3_X2 U213 ( .A1(n743), .A2(n744), .A3(in4[17]), .ZN(n1094) );
  NAND2_X2 U214 ( .A1(n549), .A2(in4[13]), .ZN(n719) );
  OAI22_X2 U215 ( .A1(n958), .A2(n959), .B1(n961), .B2(n960), .ZN(n971) );
  NAND2_X2 U216 ( .A1(n550), .A2(n551), .ZN(n575) );
  OAI211_X1 U217 ( .C1(n552), .C2(n646), .A(n619), .B(n620), .ZN(net1855) );
  INV_X4 U218 ( .A(net1861), .ZN(n552) );
  OR2_X4 U219 ( .A1(in1[28]), .A2(in3[18]), .ZN(net2879) );
  OR2_X4 U220 ( .A1(net2175), .A2(n688), .ZN(n696) );
  XOR2_X2 U221 ( .A(in1[26]), .B(in1[24]), .Z(net3004) );
  NAND3_X2 U222 ( .A1(n870), .A2(n869), .A3(in3[0]), .ZN(n679) );
  XOR2_X2 U223 ( .A(n1215), .B(n831), .Z(n1216) );
  XOR2_X2 U224 ( .A(n1203), .B(n836), .Z(n1204) );
  XOR2_X2 U225 ( .A(n1071), .B(n848), .Z(n1072) );
  XNOR2_X2 U226 ( .A(n727), .B(n762), .ZN(n1132) );
  XOR2_X1 U227 ( .A(n675), .B(n771), .Z(n1009) );
  XOR2_X1 U228 ( .A(n797), .B(n979), .Z(n980) );
  XNOR2_X1 U229 ( .A(n963), .B(n950), .ZN(n951) );
  XNOR2_X2 U230 ( .A(in4[3]), .B(n933), .ZN(n917) );
  OAI21_X2 U231 ( .B1(in4[24]), .B2(n620), .A(n644), .ZN(n553) );
  INV_X4 U232 ( .A(n553), .ZN(n637) );
  NAND2_X2 U233 ( .A1(in1[7]), .A2(in3[29]), .ZN(n739) );
  NOR2_X2 U234 ( .A1(n1076), .A2(n1077), .ZN(n746) );
  NOR2_X2 U235 ( .A1(n734), .A2(n741), .ZN(n736) );
  XNOR2_X2 U236 ( .A(in1[25]), .B(in1[27]), .ZN(n987) );
  XOR2_X2 U237 ( .A(in1[25]), .B(in1[23]), .Z(net2722) );
  XOR2_X2 U238 ( .A(n883), .B(in1[11]), .Z(n891) );
  XOR2_X2 U239 ( .A(n1186), .B(n839), .Z(n1187) );
  XOR2_X2 U240 ( .A(n1169), .B(n841), .Z(n1170) );
  XOR2_X2 U241 ( .A(n1143), .B(n843), .Z(n1144) );
  XOR2_X2 U242 ( .A(n1112), .B(n846), .Z(n1113) );
  XOR2_X2 U243 ( .A(n1090), .B(n844), .Z(n1091) );
  XOR2_X2 U244 ( .A(n1055), .B(n852), .Z(n1056) );
  OAI21_X2 U245 ( .B1(n624), .B2(n627), .A(n641), .ZN(n554) );
  INV_X4 U246 ( .A(n554), .ZN(n671) );
  XOR2_X2 U247 ( .A(n720), .B(n812), .Z(n1193) );
  AND3_X4 U248 ( .A1(n608), .A2(n606), .A3(n607), .ZN(n603) );
  XOR2_X2 U249 ( .A(n689), .B(in3[11]), .Z(net2982) );
  XNOR2_X2 U250 ( .A(in4[7]), .B(n992), .ZN(n979) );
  XNOR2_X2 U251 ( .A(n945), .B(n935), .ZN(n936) );
  XNOR2_X2 U252 ( .A(n913), .B(n899), .ZN(n900) );
  AOI211_X2 U253 ( .C1(net1722), .C2(net3978), .A(n1218), .B(n670), .ZN(
        U4_Z_30) );
  NOR2_X2 U254 ( .A1(n735), .A2(n742), .ZN(n1040) );
  NOR2_X2 U255 ( .A1(n733), .A2(n1029), .ZN(n742) );
  OR2_X4 U256 ( .A1(n596), .A2(net3065), .ZN(n555) );
  INV_X2 U257 ( .A(n1163), .ZN(n737) );
  AOI22_X1 U258 ( .A1(n985), .A2(in3[7]), .B1(n866), .B2(n833), .ZN(n865) );
  AOI21_X2 U259 ( .B1(net3479), .B2(n574), .A(n566), .ZN(net3098) );
  NAND2_X2 U260 ( .A1(n737), .A2(in4[22]), .ZN(net3421) );
  NOR2_X2 U261 ( .A1(n1028), .A2(in4[10]), .ZN(n733) );
  NOR2_X2 U262 ( .A1(n906), .A2(in3[2]), .ZN(n907) );
  OAI21_X2 U263 ( .B1(in2[28]), .B2(in4[25]), .A(net1818), .ZN(net1817) );
  AOI22_X2 U264 ( .A1(add_49_A_29_), .A2(add_49_B_29_), .B1(n1215), .B2(n591), 
        .ZN(n827) );
  AOI22_X2 U265 ( .A1(add_49_A_23_), .A2(add_49_B_23_), .B1(n1169), .B2(n581), 
        .ZN(n820) );
  AOI22_X2 U266 ( .A1(add_49_A_21_), .A2(add_49_B_21_), .B1(n1143), .B2(n577), 
        .ZN(n819) );
  AOI22_X2 U267 ( .A1(add_49_A_19_), .A2(add_49_B_19_), .B1(n1112), .B2(n576), 
        .ZN(n818) );
  OAI21_X2 U268 ( .B1(net1855), .B2(n618), .A(net1798), .ZN(n626) );
  AOI22_X2 U269 ( .A1(in1[26]), .A2(in3[16]), .B1(net3472), .B2(n807), .ZN(
        n806) );
  OAI21_X2 U270 ( .B1(n601), .B2(n602), .A(n573), .ZN(net3479) );
  NAND3_X2 U271 ( .A1(n599), .A2(n600), .A3(net3406), .ZN(n598) );
  NOR2_X2 U272 ( .A1(n701), .A2(n877), .ZN(n702) );
  INV_X4 U273 ( .A(n659), .ZN(net3979) );
  BUF_X4 U274 ( .A(n801), .Z(n711) );
  INV_X4 U275 ( .A(n779), .ZN(n1057) );
  NOR2_X2 U276 ( .A1(n1057), .A2(in4[13]), .ZN(n597) );
  AOI22_X2 U277 ( .A1(in1[8]), .A2(in3[30]), .B1(n783), .B2(n594), .ZN(n808)
         );
  INV_X4 U278 ( .A(n712), .ZN(n1019) );
  AOI22_X2 U279 ( .A1(in1[1]), .A2(in3[23]), .B1(n1158), .B2(n580), .ZN(n805)
         );
  NOR2_X2 U280 ( .A1(n710), .A2(in3[1]), .ZN(n890) );
  AOI22_X2 U281 ( .A1(add_49_A_25_), .A2(add_49_B_25_), .B1(n1186), .B2(n582), 
        .ZN(n821) );
  AOI22_X2 U282 ( .A1(add_49_A_27_), .A2(add_49_B_27_), .B1(n1203), .B2(n590), 
        .ZN(n823) );
  AOI22_X2 U283 ( .A1(add_49_A_15_), .A2(add_49_B_15_), .B1(n1071), .B2(n572), 
        .ZN(n811) );
  AOI22_X2 U284 ( .A1(add_49_A_17_), .A2(add_49_B_17_), .B1(n1090), .B2(n575), 
        .ZN(n817) );
  NOR2_X2 U285 ( .A1(n558), .A2(n559), .ZN(n556) );
  NAND2_X2 U286 ( .A1(n719), .A2(n557), .ZN(n559) );
  INV_X4 U287 ( .A(in4[14]), .ZN(n557) );
  NOR2_X2 U288 ( .A1(n559), .A2(n558), .ZN(n1064) );
  NOR2_X2 U289 ( .A1(n1058), .A2(n1059), .ZN(n558) );
  NOR2_X4 U290 ( .A1(n596), .A2(net3065), .ZN(n560) );
  INV_X1 U291 ( .A(n669), .ZN(n561) );
  INV_X4 U292 ( .A(n561), .ZN(n562) );
  AOI22_X2 U293 ( .A1(add_49_A_13_), .A2(add_49_B_13_), .B1(n1055), .B2(n571), 
        .ZN(n810) );
  NOR2_X2 U294 ( .A1(n676), .A2(in4[15]), .ZN(n1076) );
  INV_X1 U295 ( .A(n1036), .ZN(n1045) );
  AOI22_X2 U296 ( .A1(add_49_A_11_), .A2(add_49_B_11_), .B1(n1036), .B2(n569), 
        .ZN(n809) );
  INV_X1 U297 ( .A(n955), .ZN(n969) );
  AOI22_X2 U298 ( .A1(add_49_A_5_), .A2(add_49_B_5_), .B1(n955), .B2(n568), 
        .ZN(n826) );
  INV_X1 U299 ( .A(n922), .ZN(n937) );
  AOI22_X2 U300 ( .A1(add_49_A_3_), .A2(add_49_B_3_), .B1(n922), .B2(n564), 
        .ZN(n825) );
  INV_X1 U301 ( .A(n1013), .ZN(n1025) );
  AOI22_X2 U302 ( .A1(add_49_A_9_), .A2(add_49_B_9_), .B1(n1013), .B2(n570), 
        .ZN(n816) );
  INV_X4 U303 ( .A(n679), .ZN(n710) );
  INV_X1 U304 ( .A(n1158), .ZN(n1171) );
  XNOR2_X2 U305 ( .A(n966), .B(in2[9]), .ZN(n565) );
  AND2_X4 U306 ( .A1(in1[25]), .A2(in3[15]), .ZN(n566) );
  OR2_X4 U307 ( .A1(add_49_B_5_), .A2(add_49_A_5_), .ZN(n568) );
  AOI22_X2 U308 ( .A1(in1[28]), .A2(in3[18]), .B1(n567), .B2(net2879), .ZN(
        n800) );
  OR2_X4 U309 ( .A1(n605), .A2(n604), .ZN(n573) );
  OR2_X4 U310 ( .A1(in3[15]), .A2(in1[25]), .ZN(n574) );
  OR2_X4 U311 ( .A1(in3[21]), .A2(in1[31]), .ZN(n578) );
  XOR2_X2 U312 ( .A(net2175), .B(in3[10]), .Z(n579) );
  OR2_X4 U313 ( .A1(in3[23]), .A2(in1[1]), .ZN(n580) );
  AND2_X4 U314 ( .A1(n627), .A2(n641), .ZN(n583) );
  OR2_X4 U315 ( .A1(in3[26]), .A2(in1[4]), .ZN(n584) );
  XNOR2_X2 U316 ( .A(in3[30]), .B(in1[8]), .ZN(n585) );
  OR2_X4 U317 ( .A1(in4[27]), .A2(in2[30]), .ZN(n586) );
  XOR2_X2 U318 ( .A(in1[28]), .B(in3[18]), .Z(n587) );
  XOR2_X2 U319 ( .A(n605), .B(n604), .Z(n588) );
  XOR2_X2 U320 ( .A(n613), .B(n611), .Z(n589) );
  OR2_X4 U321 ( .A1(add_49_B_27_), .A2(add_49_A_27_), .ZN(n590) );
  OR2_X4 U322 ( .A1(in3[29]), .A2(in1[7]), .ZN(n592) );
  OR2_X4 U323 ( .A1(in3[27]), .A2(in1[5]), .ZN(n593) );
  OR2_X4 U324 ( .A1(in3[30]), .A2(in1[8]), .ZN(n594) );
  NOR2_X1 U325 ( .A1(n743), .A2(n744), .ZN(n595) );
  NOR2_X2 U326 ( .A1(net2882), .A2(n660), .ZN(n661) );
  AOI22_X4 U327 ( .A1(in2[30]), .A2(in4[27]), .B1(net3503), .B2(n586), .ZN(
        net2882) );
  NOR2_X2 U328 ( .A1(n1057), .A2(in4[13]), .ZN(n1058) );
  INV_X4 U329 ( .A(in3[14]), .ZN(n604) );
  XNOR2_X2 U330 ( .A(in1[24]), .B(in1[31]), .ZN(n605) );
  XNOR2_X2 U331 ( .A(n603), .B(n588), .ZN(net2094) );
  XNOR2_X2 U332 ( .A(n589), .B(n598), .ZN(net2119) );
  NAND2_X2 U333 ( .A1(n606), .A2(n607), .ZN(n601) );
  NAND2_X2 U334 ( .A1(n608), .A2(n609), .ZN(n602) );
  INV_X4 U335 ( .A(net2125), .ZN(n610) );
  INV_X4 U336 ( .A(in3[13]), .ZN(n611) );
  NAND2_X2 U337 ( .A1(n610), .A2(net4289), .ZN(n600) );
  INV_X4 U338 ( .A(n598), .ZN(n612) );
  NAND2_X2 U339 ( .A1(n613), .A2(n611), .ZN(n607) );
  NAND2_X2 U340 ( .A1(n613), .A2(n612), .ZN(n606) );
  NAND2_X2 U341 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X2 U342 ( .A1(n612), .A2(n611), .ZN(n608) );
  XNOR2_X2 U343 ( .A(in1[23]), .B(in1[30]), .ZN(n613) );
  NOR2_X1 U344 ( .A1(n874), .A2(n1210), .ZN(U5_Z_29) );
  NOR2_X2 U345 ( .A1(n631), .A2(n632), .ZN(n630) );
  NAND2_X2 U346 ( .A1(n1075), .A2(in4[15]), .ZN(n614) );
  AOI22_X2 U347 ( .A1(in1[5]), .A2(in3[27]), .B1(n724), .B2(n593), .ZN(n803)
         );
  NAND2_X2 U348 ( .A1(n614), .A2(n1084), .ZN(n731) );
  INV_X1 U349 ( .A(n895), .ZN(n615) );
  INV_X4 U350 ( .A(n615), .ZN(n616) );
  INV_X4 U351 ( .A(n894), .ZN(n895) );
  NAND3_X1 U352 ( .A1(n619), .A2(n620), .A3(n643), .ZN(n642) );
  INV_X4 U353 ( .A(n803), .ZN(n704) );
  INV_X2 U354 ( .A(n705), .ZN(n910) );
  INV_X1 U355 ( .A(n971), .ZN(n975) );
  INV_X1 U356 ( .A(n567), .ZN(n617) );
  INV_X1 U357 ( .A(n698), .ZN(net2123) );
  AND2_X2 U358 ( .A1(n808), .A2(n752), .ZN(n708) );
  NAND2_X2 U359 ( .A1(n692), .A2(n693), .ZN(net4289) );
  INV_X4 U360 ( .A(net3421), .ZN(net3196) );
  INV_X1 U361 ( .A(n691), .ZN(net3455) );
  AOI21_X4 U362 ( .B1(n621), .B2(n622), .A(n583), .ZN(net3503) );
  INV_X4 U363 ( .A(in4[24]), .ZN(n618) );
  INV_X4 U364 ( .A(net1798), .ZN(n623) );
  NOR2_X2 U365 ( .A1(n625), .A2(n626), .ZN(n624) );
  INV_X4 U366 ( .A(in4[26]), .ZN(n628) );
  NAND2_X2 U367 ( .A1(net1861), .A2(n633), .ZN(n620) );
  XNOR2_X2 U368 ( .A(in2[27]), .B(in2[31]), .ZN(n629) );
  XNOR2_X2 U369 ( .A(n629), .B(n618), .ZN(net2804) );
  XNOR2_X2 U370 ( .A(in2[16]), .B(in2[27]), .ZN(net2213) );
  XNOR2_X2 U371 ( .A(in2[17]), .B(in2[28]), .ZN(net2188) );
  XNOR2_X2 U372 ( .A(in2[29]), .B(n628), .ZN(net1815) );
  NAND2_X2 U373 ( .A1(n619), .A2(n620), .ZN(n631) );
  NAND2_X2 U374 ( .A1(n635), .A2(in4[24]), .ZN(n632) );
  NOR2_X2 U375 ( .A1(in4[24]), .A2(in4[23]), .ZN(n636) );
  NOR2_X2 U376 ( .A1(n639), .A2(n629), .ZN(n638) );
  NOR2_X2 U377 ( .A1(n623), .A2(net2902), .ZN(n622) );
  INV_X4 U378 ( .A(in4[23]), .ZN(n633) );
  NAND2_X2 U379 ( .A1(in2[29]), .A2(in4[26]), .ZN(n641) );
  INV_X4 U380 ( .A(n641), .ZN(net2902) );
  NAND2_X2 U381 ( .A1(n634), .A2(net3421), .ZN(n619) );
  NAND2_X2 U382 ( .A1(net1861), .A2(n647), .ZN(n643) );
  NAND2_X2 U383 ( .A1(net3189), .A2(net1861), .ZN(n635) );
  NAND3_X2 U384 ( .A1(net1861), .A2(net3189), .A3(n618), .ZN(n645) );
  INV_X4 U385 ( .A(n645), .ZN(n639) );
  INV_X4 U386 ( .A(n646), .ZN(n647) );
  INV_X1 U387 ( .A(net3189), .ZN(n646) );
  AOI21_X2 U388 ( .B1(n638), .B2(n637), .A(n630), .ZN(n621) );
  INV_X1 U389 ( .A(net3132), .ZN(n640) );
  NOR2_X1 U390 ( .A1(net3132), .A2(in4[23]), .ZN(n634) );
  OAI33_X1 U391 ( .A1(n662), .A2(n649), .A3(n650), .B1(n664), .B2(n651), .B3(
        n652), .ZN(n648) );
  NOR2_X2 U392 ( .A1(n648), .A2(net1690), .ZN(U4_Z_31) );
  INV_X4 U393 ( .A(n653), .ZN(n651) );
  NAND2_X2 U394 ( .A1(n665), .A2(n666), .ZN(n664) );
  OR2_X1 U395 ( .A1(net1727), .A2(n659), .ZN(n666) );
  OR2_X1 U396 ( .A1(net3065), .A2(net1727), .ZN(n667) );
  OR2_X4 U397 ( .A1(n661), .A2(n667), .ZN(n665) );
  INV_X4 U398 ( .A(n652), .ZN(n650) );
  NOR2_X2 U399 ( .A1(n650), .A2(n653), .ZN(n655) );
  OAI22_X2 U400 ( .A1(n650), .A2(net1703), .B1(n649), .B2(n655), .ZN(net1701)
         );
  INV_X4 U401 ( .A(net1703), .ZN(n649) );
  NAND2_X2 U402 ( .A1(n663), .A2(n654), .ZN(n662) );
  INV_X4 U403 ( .A(net3978), .ZN(n663) );
  XNOR2_X2 U404 ( .A(in4[31]), .B(in2[2]), .ZN(n652) );
  NAND2_X2 U405 ( .A1(n656), .A2(n657), .ZN(n653) );
  INV_X4 U406 ( .A(in4[30]), .ZN(n657) );
  INV_X4 U407 ( .A(in2[1]), .ZN(n656) );
  XOR2_X2 U408 ( .A(n656), .B(in4[30]), .Z(net1724) );
  NOR2_X2 U409 ( .A1(net1722), .A2(n659), .ZN(n658) );
  NAND2_X2 U410 ( .A1(in4[29]), .A2(in2[0]), .ZN(n654) );
  INV_X4 U411 ( .A(n654), .ZN(net1727) );
  OAI22_X2 U412 ( .A1(net1722), .A2(n654), .B1(net1727), .B2(n658), .ZN(
        net1726) );
  NOR2_X2 U413 ( .A1(in4[28]), .A2(in2[31]), .ZN(n660) );
  NOR2_X1 U414 ( .A1(n733), .A2(n1029), .ZN(n734) );
  XOR2_X2 U415 ( .A(n555), .B(n796), .Z(n1211) );
  NOR2_X2 U416 ( .A1(n560), .A2(net3979), .ZN(net3978) );
  INV_X1 U417 ( .A(net2177), .ZN(net3542) );
  NAND2_X2 U418 ( .A1(n681), .A2(n563), .ZN(n668) );
  NAND2_X2 U419 ( .A1(n681), .A2(n563), .ZN(n682) );
  NAND2_X2 U420 ( .A1(n682), .A2(n964), .ZN(n669) );
  INV_X1 U421 ( .A(net1724), .ZN(net1722) );
  INV_X4 U422 ( .A(n886), .ZN(n677) );
  NAND2_X2 U423 ( .A1(n698), .A2(in3[12]), .ZN(net3406) );
  AND2_X4 U424 ( .A1(n669), .A2(in4[6]), .ZN(n799) );
  NAND2_X2 U425 ( .A1(n702), .A2(n873), .ZN(n870) );
  INV_X4 U426 ( .A(n965), .ZN(n681) );
  INV_X1 U427 ( .A(n1075), .ZN(n672) );
  INV_X1 U428 ( .A(n999), .ZN(n673) );
  NOR2_X1 U429 ( .A1(n1004), .A2(in4[8]), .ZN(n674) );
  NOR2_X2 U430 ( .A1(n1004), .A2(in4[8]), .ZN(n1005) );
  OAI22_X2 U431 ( .A1(n678), .A2(n557), .B1(n1064), .B2(n1065), .ZN(n676) );
  NOR2_X2 U432 ( .A1(n971), .A2(in3[6]), .ZN(n972) );
  NAND2_X1 U433 ( .A1(n680), .A2(n677), .ZN(n896) );
  AND2_X4 U434 ( .A1(in4[0]), .A2(in4[1]), .ZN(n680) );
  NOR2_X4 U435 ( .A1(n963), .A2(in4[5]), .ZN(n965) );
  NAND2_X1 U436 ( .A1(n963), .A2(in4[5]), .ZN(n964) );
  NOR2_X4 U437 ( .A1(n895), .A2(in4[1]), .ZN(n897) );
  NAND2_X1 U438 ( .A1(in2[19]), .A2(n723), .ZN(n684) );
  NAND2_X2 U439 ( .A1(n683), .A2(in2[8]), .ZN(n685) );
  NAND2_X2 U440 ( .A1(n684), .A2(n685), .ZN(n792) );
  INV_X2 U441 ( .A(in2[19]), .ZN(n683) );
  INV_X2 U442 ( .A(in2[8]), .ZN(n723) );
  NAND2_X2 U443 ( .A1(n792), .A2(in2[4]), .ZN(n713) );
  INV_X2 U444 ( .A(n1004), .ZN(n1008) );
  INV_X1 U445 ( .A(n595), .ZN(n686) );
  NOR2_X2 U446 ( .A1(n1015), .A2(in3[9]), .ZN(n1016) );
  NOR2_X2 U447 ( .A1(n939), .A2(in3[4]), .ZN(n940) );
  NOR2_X4 U448 ( .A1(n945), .A2(in4[4]), .ZN(n947) );
  INV_X4 U449 ( .A(in3[10]), .ZN(n688) );
  XNOR2_X2 U450 ( .A(n690), .B(net3757), .ZN(n689) );
  XNOR2_X2 U451 ( .A(in1[21]), .B(in1[23]), .ZN(net2805) );
  XNOR2_X2 U452 ( .A(in1[21]), .B(net2489), .ZN(net2399) );
  XNOR2_X2 U453 ( .A(in1[28]), .B(in1[26]), .ZN(net2222) );
  NAND2_X2 U454 ( .A1(in3[11]), .A2(n691), .ZN(net3768) );
  INV_X4 U455 ( .A(in1[30]), .ZN(net3757) );
  NAND2_X2 U456 ( .A1(net2175), .A2(n688), .ZN(n694) );
  NAND2_X2 U457 ( .A1(net2177), .A2(n694), .ZN(n695) );
  NAND2_X2 U458 ( .A1(n695), .A2(n696), .ZN(n691) );
  NAND2_X2 U459 ( .A1(n691), .A2(n697), .ZN(n693) );
  NAND2_X2 U460 ( .A1(n697), .A2(in3[11]), .ZN(n692) );
  INV_X4 U461 ( .A(n689), .ZN(n697) );
  XNOR2_X2 U462 ( .A(in1[28]), .B(in1[21]), .ZN(n690) );
  INV_X1 U463 ( .A(n1189), .ZN(n699) );
  INV_X1 U464 ( .A(n699), .ZN(n700) );
  NAND2_X2 U465 ( .A1(n880), .A2(n879), .ZN(n786) );
  NOR2_X2 U466 ( .A1(n999), .A2(in3[8]), .ZN(n1000) );
  INV_X2 U467 ( .A(n872), .ZN(n701) );
  NAND2_X2 U468 ( .A1(n873), .A2(n872), .ZN(n703) );
  NAND2_X2 U469 ( .A1(in1[17]), .A2(in1[19]), .ZN(n872) );
  OAI22_X1 U470 ( .A1(n679), .A2(n892), .B1(n891), .B2(n890), .ZN(n705) );
  INV_X1 U471 ( .A(in1[18]), .ZN(n706) );
  NAND2_X1 U472 ( .A1(n592), .A2(n728), .ZN(n707) );
  XNOR2_X2 U473 ( .A(n804), .B(n585), .ZN(n1217) );
  NOR2_X2 U474 ( .A1(n708), .A2(n709), .ZN(U5_Z_31) );
  NAND2_X2 U475 ( .A1(n718), .A2(n876), .ZN(n709) );
  OR2_X4 U476 ( .A1(n1047), .A2(in4[12]), .ZN(n782) );
  INV_X2 U477 ( .A(n957), .ZN(n961) );
  INV_X1 U478 ( .A(in3[5]), .ZN(n960) );
  NOR2_X2 U479 ( .A1(n930), .A2(in4[3]), .ZN(n932) );
  OR2_X2 U480 ( .A1(n741), .A2(in4[11]), .ZN(n735) );
  OAI22_X1 U481 ( .A1(n673), .A2(n1002), .B1(n1000), .B2(n1001), .ZN(n712) );
  INV_X4 U482 ( .A(net3098), .ZN(net3472) );
  INV_X4 U483 ( .A(n802), .ZN(n724) );
  NAND2_X2 U484 ( .A1(n707), .A2(n739), .ZN(n714) );
  NAND2_X2 U485 ( .A1(n740), .A2(n739), .ZN(n783) );
  INV_X2 U486 ( .A(n714), .ZN(n804) );
  INV_X4 U487 ( .A(n729), .ZN(n715) );
  NAND2_X2 U488 ( .A1(n716), .A2(n717), .ZN(n718) );
  INV_X4 U489 ( .A(n808), .ZN(n716) );
  INV_X4 U490 ( .A(n752), .ZN(n717) );
  INV_X1 U491 ( .A(net2882), .ZN(net3442) );
  INV_X2 U492 ( .A(net3442), .ZN(net3443) );
  XNOR2_X2 U493 ( .A(n835), .B(in2[16]), .ZN(n1059) );
  OR2_X4 U494 ( .A1(n1022), .A2(in4[9]), .ZN(n749) );
  OAI22_X1 U495 ( .A1(n1191), .A2(n1190), .B1(n1188), .B2(n700), .ZN(n720) );
  INV_X4 U496 ( .A(n750), .ZN(n728) );
  INV_X1 U497 ( .A(n924), .ZN(n928) );
  NAND2_X1 U498 ( .A1(in2[18]), .A2(in2[7]), .ZN(n790) );
  INV_X1 U499 ( .A(n617), .ZN(n721) );
  NOR2_X2 U500 ( .A1(n726), .A2(n746), .ZN(n732) );
  INV_X2 U501 ( .A(n1160), .ZN(n1163) );
  AOI22_X2 U502 ( .A1(in1[31]), .A2(in3[21]), .B1(n1131), .B2(n578), .ZN(n801)
         );
  AOI22_X2 U503 ( .A1(in1[6]), .A2(in3[28]), .B1(n704), .B2(n751), .ZN(n750)
         );
  XOR2_X1 U504 ( .A(n1020), .B(in1[20]), .Z(net2175) );
  INV_X4 U505 ( .A(n865), .ZN(n999) );
  OR2_X2 U506 ( .A1(n985), .A2(in3[7]), .ZN(n866) );
  NAND2_X2 U507 ( .A1(n703), .A2(n877), .ZN(n869) );
  NOR2_X2 U508 ( .A1(net3196), .A2(net3132), .ZN(net3189) );
  INV_X1 U509 ( .A(n788), .ZN(n722) );
  NAND2_X2 U510 ( .A1(n728), .A2(n592), .ZN(n740) );
  XOR2_X1 U511 ( .A(n898), .B(in4[1]), .Z(n887) );
  NOR2_X2 U512 ( .A1(n913), .A2(in4[2]), .ZN(n915) );
  INV_X1 U513 ( .A(n724), .ZN(n725) );
  AOI22_X2 U514 ( .A1(in1[4]), .A2(in3[26]), .B1(n1192), .B2(n584), .ZN(n802)
         );
  INV_X1 U515 ( .A(in2[18]), .ZN(n1066) );
  INV_X2 U516 ( .A(n614), .ZN(n726) );
  OAI21_X4 U517 ( .B1(n947), .B2(n948), .A(n946), .ZN(n963) );
  OAI22_X1 U518 ( .A1(net3757), .A2(n1130), .B1(n715), .B2(n1128), .ZN(n727)
         );
  OAI22_X2 U519 ( .A1(net3757), .A2(n1130), .B1(n1129), .B2(n1128), .ZN(n1131)
         );
  NAND2_X2 U520 ( .A1(n677), .A2(in4[0]), .ZN(n894) );
  INV_X1 U521 ( .A(n1129), .ZN(n729) );
  NOR2_X2 U522 ( .A1(n1160), .A2(in4[22]), .ZN(n1161) );
  NOR2_X4 U523 ( .A1(n730), .A2(in4[7]), .ZN(n991) );
  INV_X4 U524 ( .A(n797), .ZN(n989) );
  INV_X4 U525 ( .A(n797), .ZN(n730) );
  AOI21_X4 U526 ( .B1(n798), .B2(n565), .A(n799), .ZN(n797) );
  XOR2_X1 U527 ( .A(n779), .B(n1050), .Z(n1051) );
  INV_X1 U528 ( .A(n1047), .ZN(n1049) );
  INV_X1 U529 ( .A(n737), .ZN(n738) );
  OAI21_X4 U530 ( .B1(n897), .B2(n898), .A(n896), .ZN(n913) );
  XOR2_X1 U531 ( .A(n887), .B(n616), .Z(n888) );
  OAI21_X4 U532 ( .B1(n932), .B2(n933), .A(n931), .ZN(n945) );
  NAND2_X2 U533 ( .A1(n930), .A2(in4[3]), .ZN(n931) );
  OAI21_X4 U534 ( .B1(n991), .B2(n992), .A(n990), .ZN(n1004) );
  OAI21_X4 U535 ( .B1(n915), .B2(n916), .A(n914), .ZN(n930) );
  NAND2_X2 U536 ( .A1(n913), .A2(in4[2]), .ZN(n914) );
  INV_X2 U537 ( .A(in4[10]), .ZN(n1030) );
  INV_X1 U538 ( .A(in4[16]), .ZN(n1084) );
  INV_X4 U539 ( .A(n1023), .ZN(n748) );
  INV_X1 U540 ( .A(net3479), .ZN(net2053) );
  XNOR2_X1 U541 ( .A(n647), .B(n755), .ZN(n1165) );
  INV_X1 U542 ( .A(n704), .ZN(n745) );
  AOI22_X4 U543 ( .A1(n675), .A2(in4[9]), .B1(n749), .B2(n748), .ZN(n747) );
  OR2_X1 U544 ( .A1(in3[16]), .A2(in1[26]), .ZN(n807) );
  XOR2_X2 U545 ( .A(net3004), .B(in1[17]), .Z(n833) );
  XNOR2_X2 U546 ( .A(net1855), .B(net2804), .ZN(n1174) );
  INV_X4 U547 ( .A(n753), .ZN(n824) );
  INV_X4 U548 ( .A(n754), .ZN(n828) );
  INV_X4 U549 ( .A(n757), .ZN(n822) );
  OAI22_X2 U550 ( .A1(n997), .A2(n996), .B1(n824), .B2(n995), .ZN(n757) );
  NOR2_X2 U551 ( .A1(net1750), .A2(net1751), .ZN(net3065) );
  NOR2_X2 U552 ( .A1(in3[17]), .A2(in1[27]), .ZN(n785) );
  XNOR2_X1 U553 ( .A(n721), .B(n587), .ZN(n1093) );
  OR2_X4 U554 ( .A1(in3[28]), .A2(in1[6]), .ZN(n751) );
  XNOR2_X1 U555 ( .A(n1085), .B(in2[9]), .ZN(n795) );
  XNOR2_X2 U556 ( .A(in3[31]), .B(in1[9]), .ZN(n752) );
  XNOR2_X1 U557 ( .A(in1[22]), .B(in1[24]), .ZN(n813) );
  XNOR2_X1 U558 ( .A(n1097), .B(in2[10]), .ZN(n793) );
  XNOR2_X1 U559 ( .A(net3443), .B(n814), .ZN(n1207) );
  XNOR2_X1 U560 ( .A(net1818), .B(n1181), .ZN(n1182) );
  XOR2_X1 U561 ( .A(in4[25]), .B(in2[28]), .Z(n1181) );
  OAI22_X2 U562 ( .A1(n983), .A2(n982), .B1(n826), .B2(n981), .ZN(n753) );
  OAI22_X2 U563 ( .A1(n904), .A2(n903), .B1(n902), .B2(n901), .ZN(n754) );
  XOR2_X2 U564 ( .A(in4[23]), .B(net1861), .Z(n755) );
  XNOR2_X1 U565 ( .A(n738), .B(n756), .ZN(n1153) );
  XOR2_X2 U566 ( .A(in4[22]), .B(n1162), .Z(n756) );
  XNOR2_X1 U567 ( .A(n823), .B(n832), .ZN(n1208) );
  XNOR2_X1 U568 ( .A(n1151), .B(n758), .ZN(n1139) );
  XOR2_X2 U569 ( .A(in4[21]), .B(n1149), .Z(n758) );
  XNOR2_X1 U570 ( .A(n1124), .B(n759), .ZN(n1108) );
  XOR2_X2 U571 ( .A(in4[19]), .B(n1122), .Z(n759) );
  XNOR2_X1 U572 ( .A(n1106), .B(n760), .ZN(n1098) );
  XOR2_X2 U573 ( .A(in4[18]), .B(n1104), .Z(n760) );
  XNOR2_X1 U574 ( .A(n1137), .B(n761), .ZN(n1126) );
  XOR2_X2 U575 ( .A(in4[20]), .B(n1135), .Z(n761) );
  XNOR2_X1 U576 ( .A(n834), .B(in2[15]), .ZN(n1048) );
  XNOR2_X1 U577 ( .A(n683), .B(in2[30]), .ZN(n834) );
  XNOR2_X1 U578 ( .A(n820), .B(n838), .ZN(n1175) );
  XNOR2_X1 U579 ( .A(n821), .B(n837), .ZN(n1196) );
  XOR2_X1 U580 ( .A(in3[21]), .B(in1[31]), .Z(n762) );
  XNOR2_X1 U581 ( .A(n1085), .B(in2[31]), .ZN(n835) );
  XNOR2_X1 U582 ( .A(n732), .B(n763), .ZN(n1078) );
  XOR2_X2 U583 ( .A(in4[16]), .B(n1083), .Z(n763) );
  XNOR2_X1 U584 ( .A(n687), .B(n764), .ZN(n1086) );
  XOR2_X2 U585 ( .A(in4[17]), .B(n1095), .Z(n764) );
  XOR2_X1 U586 ( .A(in3[16]), .B(in1[26]), .Z(n1073) );
  XOR2_X1 U587 ( .A(in3[17]), .B(in1[27]), .Z(n1080) );
  XNOR2_X1 U588 ( .A(n678), .B(n765), .ZN(n1060) );
  XOR2_X2 U589 ( .A(in4[14]), .B(n1065), .Z(n765) );
  XNOR2_X1 U590 ( .A(n672), .B(n766), .ZN(n1067) );
  XOR2_X2 U591 ( .A(in4[15]), .B(n1077), .Z(n766) );
  XNOR2_X1 U592 ( .A(net3542), .B(n579), .ZN(n1021) );
  XNOR2_X1 U593 ( .A(net3455), .B(net2982), .ZN(n1027) );
  XNOR2_X1 U594 ( .A(net2123), .B(n767), .ZN(n1039) );
  XOR2_X1 U595 ( .A(in3[12]), .B(net2125), .Z(n767) );
  XNOR2_X1 U596 ( .A(n736), .B(n768), .ZN(n1032) );
  XOR2_X1 U597 ( .A(in4[11]), .B(n1041), .Z(n768) );
  XNOR2_X1 U598 ( .A(n1019), .B(n769), .ZN(n1003) );
  XOR2_X1 U599 ( .A(in3[9]), .B(n1017), .Z(n769) );
  XNOR2_X1 U600 ( .A(n1008), .B(n770), .ZN(n994) );
  XOR2_X1 U601 ( .A(in4[8]), .B(n1006), .Z(n770) );
  XOR2_X1 U602 ( .A(in4[9]), .B(n1023), .Z(n771) );
  XNOR2_X1 U603 ( .A(n747), .B(n772), .ZN(n1024) );
  XOR2_X1 U604 ( .A(in4[10]), .B(n1029), .Z(n772) );
  XNOR2_X1 U605 ( .A(n673), .B(n773), .ZN(n988) );
  XOR2_X1 U606 ( .A(in3[8]), .B(n1001), .Z(n773) );
  XNOR2_X1 U607 ( .A(n975), .B(n774), .ZN(n962) );
  XOR2_X1 U608 ( .A(in3[6]), .B(n973), .Z(n774) );
  XNOR2_X1 U609 ( .A(n824), .B(n856), .ZN(n984) );
  XNOR2_X1 U610 ( .A(n822), .B(n857), .ZN(n998) );
  XNOR2_X1 U611 ( .A(n943), .B(n775), .ZN(n929) );
  XOR2_X1 U612 ( .A(in3[4]), .B(n941), .Z(n775) );
  XNOR2_X1 U613 ( .A(n961), .B(n776), .ZN(n944) );
  XOR2_X1 U614 ( .A(in3[5]), .B(n959), .Z(n776) );
  XOR2_X1 U615 ( .A(in4[5]), .B(n563), .Z(n950) );
  XNOR2_X1 U616 ( .A(n562), .B(n967), .ZN(n968) );
  XOR2_X1 U617 ( .A(in4[6]), .B(n565), .Z(n967) );
  XNOR2_X1 U618 ( .A(add_49_B_5_), .B(add_49_A_5_), .ZN(n860) );
  XNOR2_X1 U619 ( .A(n969), .B(n860), .ZN(n956) );
  XNOR2_X1 U620 ( .A(n928), .B(n777), .ZN(n912) );
  XOR2_X1 U621 ( .A(in3[3]), .B(n926), .Z(n777) );
  XNOR2_X1 U622 ( .A(n891), .B(in3[1]), .ZN(n861) );
  XOR2_X1 U623 ( .A(n861), .B(n679), .Z(n885) );
  XNOR2_X1 U624 ( .A(add_49_B_4_), .B(add_49_A_4_), .ZN(n859) );
  XNOR2_X1 U625 ( .A(n825), .B(n859), .ZN(n938) );
  XNOR2_X1 U626 ( .A(add_49_B_3_), .B(add_49_A_3_), .ZN(n858) );
  XNOR2_X1 U627 ( .A(n937), .B(n858), .ZN(n923) );
  XNOR2_X1 U628 ( .A(n910), .B(n778), .ZN(n893) );
  XOR2_X1 U629 ( .A(in3[2]), .B(n908), .Z(n778) );
  XOR2_X1 U630 ( .A(n884), .B(in3[0]), .Z(n878) );
  INV_X4 U631 ( .A(n1049), .ZN(n780) );
  INV_X4 U632 ( .A(n1048), .ZN(n781) );
  INV_X1 U633 ( .A(in1[27]), .ZN(n1092) );
  INV_X4 U634 ( .A(in3[17]), .ZN(n784) );
  AOI22_X4 U635 ( .A1(n780), .A2(in4[12]), .B1(n782), .B2(n781), .ZN(n779) );
  NAND2_X2 U636 ( .A1(n787), .A2(n786), .ZN(n886) );
  NAND2_X2 U637 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X2 U638 ( .A1(n791), .A2(n790), .ZN(n880) );
  INV_X2 U639 ( .A(in2[7]), .ZN(n788) );
  INV_X2 U640 ( .A(in2[18]), .ZN(n789) );
  INV_X4 U641 ( .A(n876), .ZN(n874) );
  INV_X4 U642 ( .A(n876), .ZN(n875) );
  XNOR2_X2 U643 ( .A(n793), .B(in2[6]), .ZN(n933) );
  XNOR2_X2 U644 ( .A(n794), .B(in1[13]), .ZN(n926) );
  XNOR2_X2 U645 ( .A(n911), .B(in1[22]), .ZN(n794) );
  XNOR2_X2 U646 ( .A(n795), .B(in2[5]), .ZN(n916) );
  XNOR2_X2 U647 ( .A(in4[29]), .B(in2[0]), .ZN(n796) );
  XNOR2_X2 U648 ( .A(in3[26]), .B(in1[4]), .ZN(n812) );
  XOR2_X2 U649 ( .A(n813), .B(in1[15]), .Z(n959) );
  XOR2_X2 U650 ( .A(net2805), .B(in1[14]), .Z(n941) );
  XNOR2_X2 U651 ( .A(in4[28]), .B(in2[31]), .ZN(n814) );
  XNOR2_X2 U652 ( .A(n671), .B(n815), .ZN(n1199) );
  XNOR2_X2 U653 ( .A(in4[27]), .B(in2[30]), .ZN(n815) );
  XNOR2_X2 U654 ( .A(n700), .B(n829), .ZN(n1180) );
  XNOR2_X2 U655 ( .A(in3[25]), .B(in1[3]), .ZN(n829) );
  XNOR2_X2 U656 ( .A(n1171), .B(n830), .ZN(n1159) );
  XNOR2_X2 U657 ( .A(in3[23]), .B(in1[1]), .ZN(n830) );
  XNOR2_X2 U658 ( .A(n987), .B(n706), .ZN(n1001) );
  XNOR2_X2 U659 ( .A(net2722), .B(in1[16]), .ZN(n973) );
  XNOR2_X2 U660 ( .A(n867), .B(n1172), .ZN(n1173) );
  XNOR2_X2 U661 ( .A(add_49_B_29_), .B(add_49_A_29_), .ZN(n831) );
  XNOR2_X2 U662 ( .A(add_49_B_28_), .B(add_49_A_28_), .ZN(n832) );
  XNOR2_X2 U663 ( .A(add_49_B_27_), .B(add_49_A_27_), .ZN(n836) );
  XNOR2_X2 U664 ( .A(add_49_B_26_), .B(add_49_A_26_), .ZN(n837) );
  XNOR2_X2 U665 ( .A(add_49_B_24_), .B(add_49_A_24_), .ZN(n838) );
  XNOR2_X2 U666 ( .A(add_49_B_25_), .B(add_49_A_25_), .ZN(n839) );
  XNOR2_X2 U667 ( .A(n819), .B(n840), .ZN(n1154) );
  XNOR2_X2 U668 ( .A(add_49_B_22_), .B(add_49_A_22_), .ZN(n840) );
  XNOR2_X2 U669 ( .A(add_49_B_23_), .B(add_49_A_23_), .ZN(n841) );
  XNOR2_X2 U670 ( .A(net2482), .B(n1073), .ZN(n1074) );
  XNOR2_X2 U671 ( .A(n868), .B(n1080), .ZN(n1081) );
  XNOR2_X2 U672 ( .A(n818), .B(n842), .ZN(n1127) );
  XNOR2_X2 U673 ( .A(add_49_B_20_), .B(add_49_A_20_), .ZN(n842) );
  XNOR2_X2 U674 ( .A(add_49_B_21_), .B(add_49_A_21_), .ZN(n843) );
  XNOR2_X2 U675 ( .A(add_49_B_17_), .B(add_49_A_17_), .ZN(n844) );
  XNOR2_X2 U676 ( .A(n817), .B(n845), .ZN(n1099) );
  XNOR2_X2 U677 ( .A(add_49_B_18_), .B(add_49_A_18_), .ZN(n845) );
  XNOR2_X2 U678 ( .A(add_49_B_19_), .B(add_49_A_19_), .ZN(n846) );
  XNOR2_X2 U679 ( .A(in4[12]), .B(n1048), .ZN(n1043) );
  XNOR2_X2 U680 ( .A(n810), .B(n847), .ZN(n1061) );
  XNOR2_X2 U681 ( .A(add_49_B_14_), .B(add_49_A_14_), .ZN(n847) );
  XNOR2_X2 U682 ( .A(add_49_B_15_), .B(add_49_A_15_), .ZN(n848) );
  XNOR2_X2 U683 ( .A(n811), .B(n849), .ZN(n1079) );
  XNOR2_X2 U684 ( .A(add_49_B_16_), .B(add_49_A_16_), .ZN(n849) );
  XNOR2_X2 U685 ( .A(in4[13]), .B(n1059), .ZN(n1050) );
  XNOR2_X2 U686 ( .A(n1045), .B(n850), .ZN(n1037) );
  XNOR2_X2 U687 ( .A(add_49_B_11_), .B(add_49_A_11_), .ZN(n850) );
  XNOR2_X2 U688 ( .A(n809), .B(n851), .ZN(n1046) );
  XNOR2_X2 U689 ( .A(add_49_B_12_), .B(add_49_A_12_), .ZN(n851) );
  XNOR2_X2 U690 ( .A(add_49_B_13_), .B(add_49_A_13_), .ZN(n852) );
  XNOR2_X2 U691 ( .A(n1025), .B(n853), .ZN(n1014) );
  XNOR2_X2 U692 ( .A(add_49_B_9_), .B(add_49_A_9_), .ZN(n853) );
  XNOR2_X2 U693 ( .A(n816), .B(n854), .ZN(n1026) );
  XNOR2_X2 U694 ( .A(add_49_B_10_), .B(add_49_A_10_), .ZN(n854) );
  XNOR2_X2 U695 ( .A(n826), .B(n855), .ZN(n970) );
  XNOR2_X2 U696 ( .A(add_49_B_6_), .B(add_49_A_6_), .ZN(n855) );
  XNOR2_X2 U697 ( .A(add_49_B_7_), .B(add_49_A_7_), .ZN(n856) );
  XNOR2_X2 U698 ( .A(add_49_B_8_), .B(add_49_A_8_), .ZN(n857) );
  AND2_X1 U699 ( .A1(n881), .A2(n876), .ZN(n862) );
  XNOR2_X2 U700 ( .A(n828), .B(n863), .ZN(n905) );
  XNOR2_X2 U701 ( .A(add_49_B_2_), .B(add_49_A_2_), .ZN(n863) );
  XOR2_X2 U702 ( .A(n864), .B(n901), .Z(n889) );
  XOR2_X2 U703 ( .A(add_49_B_1_), .B(add_49_A_1_), .Z(n864) );
  INV_X4 U704 ( .A(reset), .ZN(n876) );
  XOR2_X1 U705 ( .A(n711), .B(n1145), .Z(n1146) );
  XOR2_X1 U706 ( .A(n986), .B(n976), .Z(n977) );
  INV_X1 U707 ( .A(n985), .ZN(n986) );
  INV_X1 U708 ( .A(n939), .ZN(n943) );
  INV_X1 U709 ( .A(n1102), .ZN(n1106) );
  NOR2_X2 U710 ( .A1(n924), .A2(in3[3]), .ZN(n925) );
  INV_X1 U711 ( .A(n1120), .ZN(n1124) );
  INV_X1 U712 ( .A(n1133), .ZN(n1137) );
  INV_X1 U713 ( .A(n1147), .ZN(n1151) );
  INV_X1 U714 ( .A(n805), .ZN(n867) );
  INV_X1 U715 ( .A(net2489), .ZN(net2513) );
  INV_X2 U716 ( .A(in1[19]), .ZN(net2489) );
  INV_X1 U717 ( .A(n806), .ZN(n868) );
  INV_X1 U718 ( .A(in1[20]), .ZN(n911) );
  INV_X1 U719 ( .A(net3098), .ZN(net2482) );
  NAND2_X2 U720 ( .A1(n870), .A2(n869), .ZN(n884) );
  NAND2_X2 U721 ( .A1(n871), .A2(net2489), .ZN(n873) );
  INV_X2 U722 ( .A(in1[17]), .ZN(n871) );
  XOR2_X1 U723 ( .A(n725), .B(n1197), .Z(n1198) );
  XOR2_X1 U724 ( .A(n745), .B(n1205), .Z(n1206) );
  XOR2_X1 U725 ( .A(n750), .B(n1209), .Z(n1210) );
  XOR2_X1 U726 ( .A(net2053), .B(n1062), .Z(n1063) );
  XOR2_X1 U727 ( .A(n800), .B(n1100), .Z(n1101) );
  XOR2_X1 U728 ( .A(n715), .B(n1118), .Z(n1119) );
  INV_X4 U729 ( .A(in1[10]), .ZN(n877) );
  NOR2_X2 U730 ( .A1(n875), .A2(n878), .ZN(U5_Z_0) );
  INV_X4 U731 ( .A(in2[3]), .ZN(n879) );
  XNOR2_X2 U732 ( .A(add_49_A_0_), .B(add_49_B_0_), .ZN(n882) );
  NOR2_X2 U733 ( .A1(reset), .A2(n882), .ZN(U6_Z_0) );
  NOR2_X2 U734 ( .A1(n875), .A2(n885), .ZN(U5_Z_1) );
  NOR2_X2 U735 ( .A1(n875), .A2(n888), .ZN(U4_Z_1) );
  NAND2_X2 U736 ( .A1(add_49_B_0_), .A2(add_49_A_0_), .ZN(n901) );
  NOR2_X2 U737 ( .A1(n875), .A2(n889), .ZN(U6_Z_1) );
  INV_X4 U738 ( .A(in3[1]), .ZN(n892) );
  OAI22_X2 U739 ( .A1(n679), .A2(n892), .B1(n890), .B2(n891), .ZN(n906) );
  XNOR2_X2 U740 ( .A(net2399), .B(in1[12]), .ZN(n908) );
  NOR2_X2 U741 ( .A1(n875), .A2(n893), .ZN(U5_Z_2) );
  INV_X4 U742 ( .A(in2[20]), .ZN(n1085) );
  NOR2_X2 U743 ( .A1(n874), .A2(n900), .ZN(U4_Z_2) );
  NOR2_X2 U744 ( .A1(add_49_B_1_), .A2(add_49_A_1_), .ZN(n902) );
  NOR2_X2 U745 ( .A1(n874), .A2(n905), .ZN(U6_Z_2) );
  INV_X4 U746 ( .A(in3[2]), .ZN(n909) );
  OAI22_X2 U747 ( .A1(n910), .A2(n909), .B1(n907), .B2(n908), .ZN(n924) );
  NOR2_X2 U748 ( .A1(n875), .A2(n912), .ZN(U5_Z_3) );
  INV_X4 U749 ( .A(in2[21]), .ZN(n1097) );
  NOR2_X2 U750 ( .A1(n874), .A2(n918), .ZN(U4_Z_3) );
  NOR2_X2 U751 ( .A1(add_49_B_2_), .A2(add_49_A_2_), .ZN(n919) );
  OAI22_X2 U752 ( .A1(n921), .A2(n920), .B1(n828), .B2(n919), .ZN(n922) );
  NOR2_X2 U753 ( .A1(n875), .A2(n923), .ZN(U6_Z_3) );
  INV_X4 U754 ( .A(in3[3]), .ZN(n927) );
  OAI22_X2 U755 ( .A1(n928), .A2(n927), .B1(n925), .B2(n926), .ZN(n939) );
  NOR2_X2 U756 ( .A1(n874), .A2(n929), .ZN(U5_Z_4) );
  INV_X4 U757 ( .A(in2[22]), .ZN(n1107) );
  XOR2_X2 U758 ( .A(n1107), .B(in2[11]), .Z(n934) );
  XOR2_X2 U759 ( .A(n934), .B(n722), .Z(n948) );
  NOR2_X2 U760 ( .A1(n875), .A2(n936), .ZN(U4_Z_4) );
  NOR2_X2 U761 ( .A1(n874), .A2(n938), .ZN(U6_Z_4) );
  INV_X4 U762 ( .A(in3[4]), .ZN(n942) );
  OAI22_X2 U763 ( .A1(n943), .A2(n942), .B1(n940), .B2(n941), .ZN(n957) );
  NOR2_X2 U764 ( .A1(n875), .A2(n944), .ZN(U5_Z_5) );
  INV_X4 U765 ( .A(in2[23]), .ZN(n1125) );
  XOR2_X2 U766 ( .A(n1125), .B(in2[12]), .Z(n949) );
  NOR2_X2 U767 ( .A1(reset), .A2(n951), .ZN(U4_Z_5) );
  NOR2_X2 U768 ( .A1(add_49_B_4_), .A2(add_49_A_4_), .ZN(n952) );
  OAI22_X2 U769 ( .A1(n954), .A2(n953), .B1(n825), .B2(n952), .ZN(n955) );
  NOR2_X2 U770 ( .A1(n874), .A2(n956), .ZN(U6_Z_5) );
  NOR2_X2 U771 ( .A1(n957), .A2(in3[5]), .ZN(n958) );
  NOR2_X2 U772 ( .A1(n875), .A2(n962), .ZN(U5_Z_6) );
  INV_X4 U773 ( .A(in2[24]), .ZN(n1138) );
  XOR2_X2 U774 ( .A(n1138), .B(in2[13]), .Z(n966) );
  NOR2_X2 U775 ( .A1(n875), .A2(n968), .ZN(U4_Z_6) );
  NOR2_X2 U776 ( .A1(n874), .A2(n970), .ZN(U6_Z_6) );
  INV_X4 U777 ( .A(in3[6]), .ZN(n974) );
  OAI22_X2 U778 ( .A1(n975), .A2(n974), .B1(n972), .B2(n973), .ZN(n985) );
  XOR2_X2 U779 ( .A(in3[7]), .B(n833), .Z(n976) );
  NOR2_X2 U780 ( .A1(n875), .A2(n977), .ZN(U5_Z_7) );
  INV_X4 U781 ( .A(in2[25]), .ZN(n1152) );
  XOR2_X2 U782 ( .A(n1152), .B(in2[14]), .Z(n978) );
  XOR2_X2 U783 ( .A(n978), .B(in2[10]), .Z(n992) );
  NOR2_X2 U784 ( .A1(n874), .A2(n980), .ZN(U4_Z_7) );
  NOR2_X2 U785 ( .A1(add_49_B_6_), .A2(add_49_A_6_), .ZN(n981) );
  NOR2_X2 U786 ( .A1(n875), .A2(n984), .ZN(U6_Z_7) );
  NOR2_X2 U787 ( .A1(n875), .A2(n988), .ZN(U5_Z_8) );
  NAND2_X2 U788 ( .A1(n989), .A2(in4[7]), .ZN(n990) );
  INV_X4 U789 ( .A(in2[26]), .ZN(n1164) );
  XOR2_X2 U790 ( .A(n1164), .B(in2[15]), .Z(n993) );
  XOR2_X2 U791 ( .A(n993), .B(in2[11]), .Z(n1006) );
  NOR2_X2 U792 ( .A1(n875), .A2(n994), .ZN(U4_Z_8) );
  NOR2_X2 U793 ( .A1(add_49_B_7_), .A2(add_49_A_7_), .ZN(n995) );
  NOR2_X2 U794 ( .A1(n875), .A2(n998), .ZN(U6_Z_8) );
  INV_X4 U795 ( .A(in3[8]), .ZN(n1002) );
  OAI22_X2 U796 ( .A1(n673), .A2(n1002), .B1(n1000), .B2(n1001), .ZN(n1015) );
  XOR2_X2 U797 ( .A(net2222), .B(net2513), .Z(n1017) );
  NOR2_X2 U798 ( .A1(n875), .A2(n1003), .ZN(U5_Z_9) );
  INV_X4 U799 ( .A(in4[8]), .ZN(n1007) );
  OAI22_X2 U800 ( .A1(n1008), .A2(n1007), .B1(n1005), .B2(n1006), .ZN(n1022)
         );
  XOR2_X2 U801 ( .A(net2213), .B(in2[12]), .Z(n1023) );
  NOR2_X2 U802 ( .A1(n874), .A2(n1009), .ZN(U4_Z_9) );
  NOR2_X2 U803 ( .A1(add_49_B_8_), .A2(add_49_A_8_), .ZN(n1010) );
  OAI22_X2 U804 ( .A1(n1012), .A2(n1011), .B1(n822), .B2(n1010), .ZN(n1013) );
  NOR2_X2 U805 ( .A1(reset), .A2(n1014), .ZN(U6_Z_9) );
  INV_X4 U806 ( .A(in3[9]), .ZN(n1018) );
  OAI22_X2 U807 ( .A1(n1019), .A2(n1018), .B1(n1016), .B2(n1017), .ZN(net2177)
         );
  XOR2_X2 U808 ( .A(n1092), .B(in1[29]), .Z(n1020) );
  NOR2_X2 U809 ( .A1(n875), .A2(n1021), .ZN(U5_Z_10) );
  XOR2_X2 U810 ( .A(net2188), .B(in2[13]), .Z(n1029) );
  NOR2_X2 U811 ( .A1(reset), .A2(n1024), .ZN(U4_Z_10) );
  NOR2_X2 U812 ( .A1(n875), .A2(n1026), .ZN(U6_Z_10) );
  NOR2_X2 U813 ( .A1(n874), .A2(n1027), .ZN(U5_Z_11) );
  XOR2_X2 U814 ( .A(n1066), .B(in2[29]), .Z(n1031) );
  XOR2_X2 U815 ( .A(n1031), .B(in2[14]), .Z(n1041) );
  NOR2_X2 U816 ( .A1(n875), .A2(n1032), .ZN(U4_Z_11) );
  NOR2_X2 U817 ( .A1(add_49_B_10_), .A2(add_49_A_10_), .ZN(n1033) );
  OAI22_X2 U818 ( .A1(n1035), .A2(n1034), .B1(n816), .B2(n1033), .ZN(n1036) );
  NOR2_X2 U819 ( .A1(reset), .A2(n1037), .ZN(U6_Z_11) );
  INV_X4 U820 ( .A(in1[29]), .ZN(n1116) );
  XOR2_X2 U821 ( .A(n1116), .B(in1[31]), .Z(n1038) );
  XOR2_X2 U822 ( .A(n1038), .B(in1[22]), .Z(net2125) );
  NOR2_X2 U823 ( .A1(n874), .A2(n1039), .ZN(U5_Z_12) );
  INV_X4 U824 ( .A(in4[11]), .ZN(n1042) );
  OAI22_X2 U825 ( .A1(n736), .A2(n1042), .B1(n1040), .B2(n1041), .ZN(n1047) );
  XOR2_X2 U826 ( .A(n1049), .B(n1043), .Z(n1044) );
  NOR2_X2 U827 ( .A1(n875), .A2(n1044), .ZN(U4_Z_12) );
  NOR2_X2 U828 ( .A1(n874), .A2(n1046), .ZN(U6_Z_12) );
  NOR2_X2 U829 ( .A1(n875), .A2(net2119), .ZN(U5_Z_13) );
  NOR2_X2 U830 ( .A1(n875), .A2(n1051), .ZN(U4_Z_13) );
  NOR2_X2 U831 ( .A1(add_49_B_12_), .A2(add_49_A_12_), .ZN(n1052) );
  OAI22_X2 U832 ( .A1(n1054), .A2(n1053), .B1(n809), .B2(n1052), .ZN(n1055) );
  NOR2_X2 U833 ( .A1(n874), .A2(n1056), .ZN(U6_Z_13) );
  NOR2_X2 U834 ( .A1(n875), .A2(net2094), .ZN(U5_Z_14) );
  XOR2_X2 U835 ( .A(n1097), .B(in2[17]), .Z(n1065) );
  NOR2_X2 U836 ( .A1(n875), .A2(n1060), .ZN(U4_Z_14) );
  NOR2_X2 U837 ( .A1(n874), .A2(n1061), .ZN(U6_Z_14) );
  XOR2_X2 U838 ( .A(in3[15]), .B(in1[25]), .Z(n1062) );
  NOR2_X2 U839 ( .A1(n875), .A2(n1063), .ZN(U5_Z_15) );
  OAI22_X2 U840 ( .A1(n678), .A2(n557), .B1(n556), .B2(n1065), .ZN(n1075) );
  XOR2_X2 U841 ( .A(n1066), .B(in2[22]), .Z(n1077) );
  NOR2_X2 U842 ( .A1(n875), .A2(n1067), .ZN(U4_Z_15) );
  NOR2_X2 U843 ( .A1(add_49_B_14_), .A2(add_49_A_14_), .ZN(n1068) );
  OAI22_X2 U844 ( .A1(n1070), .A2(n1069), .B1(n810), .B2(n1068), .ZN(n1071) );
  NOR2_X2 U845 ( .A1(n875), .A2(n1072), .ZN(U6_Z_15) );
  NOR2_X2 U846 ( .A1(n874), .A2(n1074), .ZN(U5_Z_16) );
  XOR2_X2 U847 ( .A(n683), .B(in2[23]), .Z(n1083) );
  NOR2_X2 U848 ( .A1(n874), .A2(n1078), .ZN(U4_Z_16) );
  NOR2_X2 U849 ( .A1(n874), .A2(n1079), .ZN(U6_Z_16) );
  NOR2_X2 U850 ( .A1(n874), .A2(n1081), .ZN(U5_Z_17) );
  NOR2_X2 U851 ( .A1(n746), .A2(n731), .ZN(n1082) );
  XOR2_X2 U852 ( .A(n1085), .B(in2[24]), .Z(n1095) );
  NOR2_X2 U853 ( .A1(n874), .A2(n1086), .ZN(U4_Z_17) );
  NOR2_X2 U854 ( .A1(add_49_B_16_), .A2(add_49_A_16_), .ZN(n1087) );
  OAI22_X2 U855 ( .A1(n1089), .A2(n1088), .B1(n811), .B2(n1087), .ZN(n1090) );
  NOR2_X2 U856 ( .A1(n874), .A2(n1091), .ZN(U6_Z_17) );
  NOR2_X2 U857 ( .A1(n874), .A2(n1093), .ZN(U5_Z_18) );
  INV_X4 U858 ( .A(in4[17]), .ZN(n1096) );
  OAI22_X2 U859 ( .A1(n687), .A2(n1096), .B1(n1094), .B2(n1095), .ZN(n1102) );
  XOR2_X2 U860 ( .A(n1097), .B(in2[25]), .Z(n1104) );
  NOR2_X2 U861 ( .A1(n874), .A2(n1098), .ZN(U4_Z_18) );
  NOR2_X2 U862 ( .A1(n874), .A2(n1099), .ZN(U6_Z_18) );
  XOR2_X2 U863 ( .A(in3[19]), .B(in1[29]), .Z(n1100) );
  NOR2_X2 U864 ( .A1(n874), .A2(n1101), .ZN(U5_Z_19) );
  INV_X4 U865 ( .A(in4[18]), .ZN(n1105) );
  NOR2_X2 U866 ( .A1(n1102), .A2(in4[18]), .ZN(n1103) );
  OAI22_X2 U867 ( .A1(n1106), .A2(n1105), .B1(n1103), .B2(n1104), .ZN(n1120)
         );
  XOR2_X2 U868 ( .A(n1107), .B(in2[26]), .Z(n1122) );
  NOR2_X2 U869 ( .A1(n874), .A2(n1108), .ZN(U4_Z_19) );
  NOR2_X2 U870 ( .A1(add_49_B_18_), .A2(add_49_A_18_), .ZN(n1109) );
  OAI22_X2 U871 ( .A1(n1111), .A2(n1110), .B1(n817), .B2(n1109), .ZN(n1112) );
  NOR2_X2 U872 ( .A1(n874), .A2(n1113), .ZN(U6_Z_19) );
  INV_X4 U873 ( .A(in3[19]), .ZN(n1115) );
  NOR2_X2 U874 ( .A1(in3[19]), .A2(in1[29]), .ZN(n1114) );
  OAI22_X2 U875 ( .A1(n1116), .A2(n1115), .B1(n800), .B2(n1114), .ZN(n1117) );
  INV_X4 U876 ( .A(n1117), .ZN(n1129) );
  XOR2_X2 U877 ( .A(in3[20]), .B(in1[30]), .Z(n1118) );
  NOR2_X2 U878 ( .A1(n874), .A2(n1119), .ZN(U5_Z_20) );
  INV_X4 U879 ( .A(in4[19]), .ZN(n1123) );
  NOR2_X2 U880 ( .A1(n1120), .A2(in4[19]), .ZN(n1121) );
  OAI22_X2 U881 ( .A1(n1124), .A2(n1123), .B1(n1121), .B2(n1122), .ZN(n1133)
         );
  XOR2_X2 U882 ( .A(n1125), .B(in2[27]), .Z(n1135) );
  NOR2_X2 U883 ( .A1(n874), .A2(n1126), .ZN(U4_Z_20) );
  NOR2_X2 U884 ( .A1(n874), .A2(n1127), .ZN(U6_Z_20) );
  INV_X4 U885 ( .A(in3[20]), .ZN(n1130) );
  NOR2_X2 U886 ( .A1(in3[20]), .A2(in1[30]), .ZN(n1128) );
  NOR2_X2 U887 ( .A1(n875), .A2(n1132), .ZN(U5_Z_21) );
  INV_X4 U888 ( .A(in4[20]), .ZN(n1136) );
  NOR2_X2 U889 ( .A1(n1133), .A2(in4[20]), .ZN(n1134) );
  OAI22_X2 U890 ( .A1(n1137), .A2(n1136), .B1(n1134), .B2(n1135), .ZN(n1147)
         );
  XOR2_X2 U891 ( .A(n1138), .B(in2[28]), .Z(n1149) );
  NOR2_X2 U892 ( .A1(n874), .A2(n1139), .ZN(U4_Z_21) );
  NOR2_X2 U893 ( .A1(add_49_B_20_), .A2(add_49_A_20_), .ZN(n1140) );
  OAI22_X2 U894 ( .A1(n1142), .A2(n1141), .B1(n818), .B2(n1140), .ZN(n1143) );
  NOR2_X2 U895 ( .A1(reset), .A2(n1144), .ZN(U6_Z_21) );
  XOR2_X2 U896 ( .A(in3[22]), .B(in1[0]), .Z(n1145) );
  NOR2_X2 U897 ( .A1(n874), .A2(n1146), .ZN(U5_Z_22) );
  INV_X4 U898 ( .A(in4[21]), .ZN(n1150) );
  NOR2_X2 U899 ( .A1(n1147), .A2(in4[21]), .ZN(n1148) );
  OAI22_X2 U900 ( .A1(n1151), .A2(n1150), .B1(n1148), .B2(n1149), .ZN(n1160)
         );
  XOR2_X2 U901 ( .A(n1152), .B(in2[29]), .Z(n1162) );
  NOR2_X2 U902 ( .A1(n874), .A2(n1153), .ZN(U4_Z_22) );
  NOR2_X2 U903 ( .A1(n874), .A2(n1154), .ZN(U6_Z_22) );
  INV_X4 U904 ( .A(in1[0]), .ZN(n1157) );
  INV_X4 U905 ( .A(in3[22]), .ZN(n1156) );
  NOR2_X2 U906 ( .A1(in3[22]), .A2(in1[0]), .ZN(n1155) );
  OAI22_X2 U907 ( .A1(n1157), .A2(n1156), .B1(n801), .B2(n1155), .ZN(n1158) );
  NOR2_X2 U908 ( .A1(n875), .A2(n1159), .ZN(U5_Z_23) );
  XOR2_X2 U909 ( .A(n1164), .B(in2[30]), .Z(net1861) );
  NOR2_X2 U910 ( .A1(reset), .A2(n1165), .ZN(U4_Z_23) );
  NOR2_X2 U911 ( .A1(add_49_B_22_), .A2(add_49_A_22_), .ZN(n1166) );
  OAI22_X2 U912 ( .A1(n1168), .A2(n1167), .B1(n819), .B2(n1166), .ZN(n1169) );
  NOR2_X2 U913 ( .A1(n874), .A2(n1170), .ZN(U6_Z_23) );
  XOR2_X2 U914 ( .A(in3[24]), .B(in1[2]), .Z(n1172) );
  NOR2_X2 U915 ( .A1(reset), .A2(n1173), .ZN(U5_Z_24) );
  NOR2_X2 U916 ( .A1(n874), .A2(n1174), .ZN(U4_Z_24) );
  NOR2_X2 U917 ( .A1(n874), .A2(n1175), .ZN(U6_Z_24) );
  INV_X4 U918 ( .A(in1[2]), .ZN(n1178) );
  INV_X4 U919 ( .A(in3[24]), .ZN(n1177) );
  NOR2_X2 U920 ( .A1(in3[24]), .A2(in1[2]), .ZN(n1176) );
  OAI22_X2 U921 ( .A1(n1178), .A2(n1177), .B1(n805), .B2(n1176), .ZN(n1179) );
  INV_X4 U922 ( .A(n1179), .ZN(n1189) );
  NOR2_X2 U923 ( .A1(n874), .A2(n1180), .ZN(U5_Z_25) );
  NOR2_X2 U924 ( .A1(n874), .A2(n1182), .ZN(U4_Z_25) );
  NOR2_X2 U925 ( .A1(add_49_B_24_), .A2(add_49_A_24_), .ZN(n1183) );
  OAI22_X2 U926 ( .A1(n1185), .A2(n1184), .B1(n820), .B2(n1183), .ZN(n1186) );
  NOR2_X2 U927 ( .A1(n874), .A2(n1187), .ZN(U6_Z_25) );
  INV_X4 U928 ( .A(in1[3]), .ZN(n1191) );
  INV_X4 U929 ( .A(in3[25]), .ZN(n1190) );
  NOR2_X2 U930 ( .A1(in3[25]), .A2(in1[3]), .ZN(n1188) );
  OAI22_X2 U931 ( .A1(n1191), .A2(n1190), .B1(n1189), .B2(n1188), .ZN(n1192)
         );
  NOR2_X2 U932 ( .A1(n874), .A2(n1193), .ZN(U5_Z_26) );
  NAND2_X2 U933 ( .A1(in4[25]), .A2(in2[28]), .ZN(net1798) );
  NAND2_X2 U934 ( .A1(net1798), .A2(net1817), .ZN(n1194) );
  XNOR2_X2 U935 ( .A(net1815), .B(n1194), .ZN(n1195) );
  NOR2_X2 U936 ( .A1(n874), .A2(n1195), .ZN(U4_Z_26) );
  NOR2_X2 U937 ( .A1(n874), .A2(n1196), .ZN(U6_Z_26) );
  XOR2_X2 U938 ( .A(in3[27]), .B(in1[5]), .Z(n1197) );
  NOR2_X2 U939 ( .A1(n874), .A2(n1198), .ZN(U5_Z_27) );
  NOR2_X2 U940 ( .A1(n874), .A2(n1199), .ZN(U4_Z_27) );
  NOR2_X2 U941 ( .A1(add_49_B_26_), .A2(add_49_A_26_), .ZN(n1200) );
  OAI22_X2 U942 ( .A1(n1202), .A2(n1201), .B1(n821), .B2(n1200), .ZN(n1203) );
  NOR2_X2 U943 ( .A1(n874), .A2(n1204), .ZN(U6_Z_27) );
  XOR2_X2 U944 ( .A(in3[28]), .B(in1[6]), .Z(n1205) );
  NOR2_X2 U945 ( .A1(n874), .A2(n1206), .ZN(U5_Z_28) );
  NOR2_X2 U946 ( .A1(n875), .A2(n1207), .ZN(U4_Z_28) );
  NOR2_X2 U947 ( .A1(n875), .A2(n1208), .ZN(U6_Z_28) );
  XOR2_X2 U948 ( .A(in3[29]), .B(in1[7]), .Z(n1209) );
  INV_X4 U949 ( .A(in2[31]), .ZN(net1750) );
  INV_X4 U950 ( .A(in4[28]), .ZN(net1751) );
  NOR2_X2 U951 ( .A1(reset), .A2(n1211), .ZN(U4_Z_29) );
  NOR2_X2 U952 ( .A1(add_49_B_28_), .A2(add_49_A_28_), .ZN(n1212) );
  OAI22_X2 U953 ( .A1(n1214), .A2(n1213), .B1(n823), .B2(n1212), .ZN(n1215) );
  NOR2_X2 U954 ( .A1(reset), .A2(n1216), .ZN(U6_Z_29) );
  NOR2_X2 U955 ( .A1(n874), .A2(n1217), .ZN(U5_Z_30) );
  NAND2_X2 U956 ( .A1(net1726), .A2(n876), .ZN(n1218) );
  XOR2_X2 U957 ( .A(add_49_B_30_), .B(add_49_A_30_), .Z(n1219) );
  XOR2_X2 U958 ( .A(n827), .B(n1219), .Z(n1220) );
  NOR2_X2 U959 ( .A1(reset), .A2(n1220), .ZN(U6_Z_30) );
  NAND2_X2 U960 ( .A1(in4[30]), .A2(in2[1]), .ZN(net1703) );
  NAND2_X2 U961 ( .A1(net1701), .A2(n876), .ZN(net1690) );
  XNOR2_X2 U962 ( .A(add_49_B_31_), .B(add_49_A_31_), .ZN(n1225) );
  NOR2_X2 U963 ( .A1(add_49_B_30_), .A2(add_49_A_30_), .ZN(n1221) );
  OAI22_X2 U964 ( .A1(n1223), .A2(n1222), .B1(n827), .B2(n1221), .ZN(n1224) );
  XOR2_X2 U965 ( .A(n1225), .B(n1224), .Z(n1226) );
  NOR2_X2 U966 ( .A1(reset), .A2(n1226), .ZN(U6_Z_31) );
endmodule

