
module fp_1 ( clock, reset, in1, in2, in3, in4, ops_out );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  output [31:0] ops_out;
  input clock, reset;
  wire   U9_Z_0, U9_Z_1, U9_Z_2, U9_Z_3, U9_Z_4, U9_Z_5, U9_Z_6, U9_Z_7,
         U9_Z_8, U9_Z_9, U9_Z_10, U9_Z_11, U9_Z_12, U9_Z_13, U9_Z_14, U9_Z_15,
         U9_Z_16, U9_Z_17, U9_Z_18, U9_Z_19, U9_Z_20, U9_Z_21, U9_Z_22,
         U9_Z_23, U9_Z_24, U9_Z_25, U9_Z_26, U9_Z_27, U9_Z_28, U9_Z_29,
         U9_Z_30, U9_Z_31, U8_Z_0, U8_Z_1, U8_Z_2, U8_Z_3, U8_Z_4, U8_Z_5,
         U8_Z_6, U8_Z_7, U8_Z_8, U8_Z_9, U8_Z_10, U8_Z_11, U8_Z_12, U8_Z_13,
         U8_Z_14, U8_Z_15, U8_Z_16, U8_Z_17, U8_Z_18, U8_Z_19, U8_Z_20,
         U8_Z_21, U8_Z_22, U8_Z_23, U8_Z_24, U8_Z_25, U8_Z_26, U8_Z_27,
         U8_Z_28, U8_Z_29, U8_Z_30, U8_Z_31, U7_Z_1, U7_Z_2, U7_Z_3, U7_Z_4,
         U7_Z_5, U7_Z_6, U7_Z_7, U7_Z_8, U7_Z_9, U7_Z_10, U7_Z_11, U7_Z_12,
         U7_Z_13, U7_Z_14, U7_Z_15, U7_Z_16, U7_Z_17, U7_Z_18, U7_Z_19,
         U7_Z_20, U7_Z_21, U7_Z_22, U7_Z_23, U7_Z_24, U7_Z_25, U7_Z_26,
         U7_Z_27, U7_Z_28, U7_Z_29, U7_Z_30, U7_Z_31, U6_A_31_, U6_A_30_,
         U6_A_29_, U6_A_28_, U6_A_27_, U6_A_26_, U6_A_25_, U6_A_24_, U6_A_23_,
         U6_A_22_, U6_A_21_, U6_A_20_, U6_A_19_, U6_A_18_, U6_A_17_, U6_A_16_,
         U6_A_15_, U6_A_14_, U6_A_13_, U6_A_12_, U6_A_11_, U6_A_10_, U6_A_9_,
         U6_A_8_, U6_A_7_, U6_A_6_, U6_A_5_, U6_A_4_, U6_A_3_, U6_A_2_,
         U6_A_1_, U6_A_0_, U6_B_31_, U6_B_30_, U6_B_29_, U6_B_28_, U6_B_27_,
         U6_B_26_, U6_B_25_, U6_B_24_, U6_B_23_, U6_B_22_, U6_B_21_, U6_B_20_,
         U6_B_19_, U6_B_18_, U6_B_17_, U6_B_16_, U6_B_15_, U6_B_14_, U6_B_13_,
         U6_B_12_, U6_B_11_, U6_B_10_, U6_B_9_, U6_B_8_, U6_B_7_, U6_B_6_,
         U6_B_5_, U6_B_4_, U6_B_3_, U6_B_2_, U6_B_1_, U6_B_0_, net3512,
         net3523, net3525, net3544, net3546, net3548, net3549, net3572,
         net3573, net3620, net3637, net3639, net3640, net3677, net3683,
         net3875, net3916, net3941, net3945, net3947, net3997, net3999,
         net4010, net4035, net4044, net4221, net4311, net4304, net4335,
         net4544, net4626, net4627, net4701, net4704, net4724, net4804,
         net4826, net4887, net4920, net4954, net5011, net5018, net5228,
         net5243, net5265, net5264, net5277, net5294, net5301, net5325,
         net5364, net5590, net5579, net5801, net5800, net6111, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325;

  DFF_X2 adr_2_op_reg_30_ ( .D(U7_Z_30), .CK(clock), .Q(U6_B_30_), .QN(n1321)
         );
  DFF_X2 adr_2_op_reg_0_ ( .D(n961), .CK(clock), .Q(U6_B_0_) );
  DFF_X2 adr_1_op_reg_0_ ( .D(U8_Z_0), .CK(clock), .Q(U6_A_0_) );
  DFF_X2 adr_1_op_reg_1_ ( .D(U8_Z_1), .CK(clock), .Q(U6_A_1_), .QN(n1003) );
  DFF_X2 adr_2_op_reg_3_ ( .D(U7_Z_3), .CK(clock), .Q(U6_B_3_), .QN(n637) );
  DFF_X2 adr_2_op_reg_2_ ( .D(U7_Z_2), .CK(clock), .Q(U6_B_2_), .QN(n1019) );
  DFF_X2 adr_2_op_reg_1_ ( .D(U7_Z_1), .CK(clock), .Q(U6_B_1_), .QN(n1002) );
  DFF_X2 adr_1_op_reg_2_ ( .D(U8_Z_2), .CK(clock), .Q(U6_A_2_), .QN(n1020) );
  DFF_X2 adr_2_op_reg_4_ ( .D(U7_Z_4), .CK(clock), .Q(U6_B_4_), .QN(n1052) );
  DFF_X2 adr_1_op_reg_3_ ( .D(U8_Z_3), .CK(clock), .Q(U6_A_3_), .QN(n638) );
  DFF_X2 adr_2_op_reg_5_ ( .D(U7_Z_5), .CK(clock), .Q(U6_B_5_) );
  DFF_X2 adr_1_op_reg_4_ ( .D(U8_Z_4), .CK(clock), .Q(U6_A_4_), .QN(n1053) );
  DFF_X2 adr_1_op_reg_5_ ( .D(U8_Z_5), .CK(clock), .Q(U6_A_5_) );
  DFF_X2 adr_2_op_reg_7_ ( .D(U7_Z_7), .CK(clock), .Q(U6_B_7_), .QN(n1095) );
  DFF_X2 adr_2_op_reg_6_ ( .D(U7_Z_6), .CK(clock), .Q(U6_B_6_), .QN(n1081) );
  DFF_X2 adr_2_op_reg_8_ ( .D(U7_Z_8), .CK(clock), .Q(U6_B_8_), .QN(n1110) );
  DFF_X2 adr_1_op_reg_6_ ( .D(U8_Z_6), .CK(clock), .Q(U6_A_6_), .QN(n1082) );
  DFF_X2 adr_2_op_reg_9_ ( .D(U7_Z_9), .CK(clock), .Q(U6_B_9_), .QN(n635) );
  DFF_X2 adr_1_op_reg_7_ ( .D(U8_Z_7), .CK(clock), .Q(U6_A_7_), .QN(n1096) );
  DFF_X2 adr_1_op_reg_8_ ( .D(U8_Z_8), .CK(clock), .Q(U6_A_8_), .QN(n1111) );
  DFF_X2 adr_2_op_reg_10_ ( .D(U7_Z_10), .CK(clock), .Q(U6_B_10_), .QN(n1133)
         );
  DFF_X2 adr_2_op_reg_11_ ( .D(U7_Z_11), .CK(clock), .Q(U6_B_11_), .QN(n645)
         );
  DFF_X2 adr_1_op_reg_10_ ( .D(U8_Z_10), .CK(clock), .Q(U6_A_10_), .QN(n1134)
         );
  DFF_X2 adr_1_op_reg_9_ ( .D(U8_Z_9), .CK(clock), .Q(U6_A_9_), .QN(n636) );
  DFF_X2 adr_2_op_reg_12_ ( .D(U7_Z_12), .CK(clock), .Q(U6_B_12_), .QN(n1152)
         );
  DFF_X2 adr_1_op_reg_11_ ( .D(U8_Z_11), .CK(clock), .Q(U6_A_11_), .QN(n646)
         );
  DFF_X2 adr_1_op_reg_12_ ( .D(U8_Z_12), .CK(clock), .Q(U6_A_12_), .QN(n1153)
         );
  DFF_X2 adr_1_op_reg_13_ ( .D(U8_Z_13), .CK(clock), .Q(U6_A_13_), .QN(n629)
         );
  DFF_X2 adr_2_op_reg_13_ ( .D(U7_Z_13), .CK(clock), .Q(U6_B_13_), .QN(n628)
         );
  DFF_X2 adr_2_op_reg_14_ ( .D(U7_Z_14), .CK(clock), .Q(U6_B_14_), .QN(n1168)
         );
  DFF_X2 adr_1_op_reg_14_ ( .D(U8_Z_14), .CK(clock), .Q(U6_A_14_), .QN(n1169)
         );
  DFF_X2 adr_1_op_reg_15_ ( .D(U8_Z_15), .CK(clock), .Q(U6_A_15_), .QN(n634)
         );
  DFF_X2 adr_1_op_reg_16_ ( .D(U8_Z_16), .CK(clock), .Q(U6_A_16_), .QN(n1188)
         );
  DFF_X2 adr_2_op_reg_15_ ( .D(U7_Z_15), .CK(clock), .Q(U6_B_15_), .QN(n633)
         );
  DFF_X2 adr_1_op_reg_17_ ( .D(U8_Z_17), .CK(clock), .Q(U6_A_17_), .QN(n650)
         );
  DFF_X2 adr_2_op_reg_16_ ( .D(U7_Z_16), .CK(clock), .Q(U6_B_16_), .QN(n1187)
         );
  DFF_X2 adr_1_op_reg_18_ ( .D(U8_Z_18), .CK(clock), .Q(U6_A_18_), .QN(n1210)
         );
  DFF_X2 adr_2_op_reg_17_ ( .D(U7_Z_17), .CK(clock), .Q(U6_B_17_), .QN(n649)
         );
  DFF_X2 adr_1_op_reg_19_ ( .D(U8_Z_19), .CK(clock), .Q(U6_A_19_), .QN(n644)
         );
  DFF_X2 adr_2_op_reg_18_ ( .D(U7_Z_18), .CK(clock), .Q(U6_B_18_), .QN(n1209)
         );
  DFF_X2 adr_1_op_reg_20_ ( .D(U8_Z_20), .CK(clock), .Q(U6_A_20_), .QN(n1241)
         );
  DFF_X2 adr_2_op_reg_19_ ( .D(U7_Z_19), .CK(clock), .Q(U6_B_19_), .QN(n643)
         );
  DFF_X2 adr_2_op_reg_20_ ( .D(U7_Z_20), .CK(clock), .Q(U6_B_20_), .QN(n1240)
         );
  DFF_X2 adr_1_op_reg_21_ ( .D(U8_Z_21), .CK(clock), .Q(U6_A_21_), .QN(n632)
         );
  DFF_X2 adr_2_op_reg_21_ ( .D(U7_Z_21), .CK(clock), .Q(U6_B_21_), .QN(n631)
         );
  DFF_X2 adr_1_op_reg_22_ ( .D(U8_Z_22), .CK(clock), .Q(U6_A_22_), .QN(n1267)
         );
  DFF_X2 adr_1_op_reg_23_ ( .D(U8_Z_23), .CK(clock), .Q(U6_A_23_), .QN(n627)
         );
  DFF_X2 adr_2_op_reg_22_ ( .D(U7_Z_22), .CK(clock), .Q(U6_B_22_), .QN(n1266)
         );
  DFF_X2 adr_1_op_reg_24_ ( .D(U8_Z_24), .CK(clock), .Q(U6_A_24_), .QN(n1284)
         );
  DFF_X2 adr_2_op_reg_23_ ( .D(U7_Z_23), .CK(clock), .Q(U6_B_23_), .QN(n626)
         );
  DFF_X2 adr_1_op_reg_25_ ( .D(U8_Z_25), .CK(clock), .Q(U6_A_25_), .QN(n642)
         );
  DFF_X2 adr_2_op_reg_24_ ( .D(U7_Z_24), .CK(clock), .Q(U6_B_24_), .QN(n1283)
         );
  DFF_X2 adr_1_op_reg_27_ ( .D(U8_Z_27), .CK(clock), .Q(U6_A_27_) );
  DFF_X2 adr_1_op_reg_26_ ( .D(U8_Z_26), .CK(clock), .Q(U6_A_26_), .QN(n1301)
         );
  DFF_X2 adr_1_op_reg_28_ ( .D(U8_Z_28), .CK(clock), .Q(U6_A_28_), .QN(n1313)
         );
  DFF_X2 adr_2_op_reg_27_ ( .D(U7_Z_27), .CK(clock), .Q(U6_B_27_) );
  DFF_X2 adr_1_op_reg_29_ ( .D(U8_Z_29), .CK(clock), .Q(U6_A_29_), .QN(n625)
         );
  DFF_X2 adr_1_op_reg_30_ ( .D(U8_Z_30), .CK(clock), .Q(U6_A_30_), .QN(n1322)
         );
  DFF_X2 adr_2_op_reg_28_ ( .D(U7_Z_28), .CK(clock), .Q(U6_B_28_), .QN(n1312)
         );
  DFF_X2 adr_2_op_reg_29_ ( .D(U7_Z_29), .CK(clock), .Q(U6_B_29_), .QN(n624)
         );
  DFF_X2 ops_out_reg_0_ ( .D(U9_Z_0), .CK(clock), .Q(ops_out[0]) );
  DFF_X2 ops_out_reg_2_ ( .D(U9_Z_2), .CK(clock), .Q(ops_out[2]) );
  DFF_X2 ops_out_reg_1_ ( .D(U9_Z_1), .CK(clock), .Q(ops_out[1]) );
  DFF_X2 ops_out_reg_3_ ( .D(U9_Z_3), .CK(clock), .Q(ops_out[3]) );
  DFF_X2 ops_out_reg_4_ ( .D(U9_Z_4), .CK(clock), .Q(ops_out[4]) );
  DFF_X2 ops_out_reg_5_ ( .D(U9_Z_5), .CK(clock), .Q(ops_out[5]) );
  DFF_X2 ops_out_reg_6_ ( .D(U9_Z_6), .CK(clock), .Q(ops_out[6]) );
  DFF_X2 ops_out_reg_7_ ( .D(U9_Z_7), .CK(clock), .Q(ops_out[7]) );
  DFF_X2 ops_out_reg_8_ ( .D(U9_Z_8), .CK(clock), .Q(ops_out[8]) );
  DFF_X2 ops_out_reg_9_ ( .D(U9_Z_9), .CK(clock), .Q(ops_out[9]) );
  DFF_X2 ops_out_reg_10_ ( .D(U9_Z_10), .CK(clock), .Q(ops_out[10]) );
  DFF_X2 ops_out_reg_11_ ( .D(U9_Z_11), .CK(clock), .Q(ops_out[11]) );
  DFF_X2 ops_out_reg_12_ ( .D(U9_Z_12), .CK(clock), .Q(ops_out[12]) );
  DFF_X2 ops_out_reg_13_ ( .D(U9_Z_13), .CK(clock), .Q(ops_out[13]) );
  DFF_X2 ops_out_reg_14_ ( .D(U9_Z_14), .CK(clock), .Q(ops_out[14]) );
  DFF_X2 ops_out_reg_15_ ( .D(U9_Z_15), .CK(clock), .Q(ops_out[15]) );
  DFF_X2 ops_out_reg_16_ ( .D(U9_Z_16), .CK(clock), .Q(ops_out[16]) );
  DFF_X2 ops_out_reg_17_ ( .D(U9_Z_17), .CK(clock), .Q(ops_out[17]) );
  DFF_X2 ops_out_reg_18_ ( .D(U9_Z_18), .CK(clock), .Q(ops_out[18]) );
  DFF_X2 ops_out_reg_19_ ( .D(U9_Z_19), .CK(clock), .Q(ops_out[19]) );
  DFF_X2 ops_out_reg_20_ ( .D(U9_Z_20), .CK(clock), .Q(ops_out[20]) );
  DFF_X2 ops_out_reg_21_ ( .D(U9_Z_21), .CK(clock), .Q(ops_out[21]) );
  DFF_X2 ops_out_reg_22_ ( .D(U9_Z_22), .CK(clock), .Q(ops_out[22]) );
  DFF_X2 ops_out_reg_23_ ( .D(U9_Z_23), .CK(clock), .Q(ops_out[23]) );
  DFF_X2 ops_out_reg_24_ ( .D(U9_Z_24), .CK(clock), .Q(ops_out[24]) );
  DFF_X2 ops_out_reg_25_ ( .D(U9_Z_25), .CK(clock), .Q(ops_out[25]) );
  DFF_X2 ops_out_reg_26_ ( .D(U9_Z_26), .CK(clock), .Q(ops_out[26]) );
  DFF_X2 ops_out_reg_27_ ( .D(U9_Z_27), .CK(clock), .Q(ops_out[27]) );
  DFF_X2 ops_out_reg_28_ ( .D(U9_Z_28), .CK(clock), .Q(ops_out[28]) );
  DFF_X2 ops_out_reg_29_ ( .D(U9_Z_29), .CK(clock), .Q(ops_out[29]) );
  DFF_X2 ops_out_reg_30_ ( .D(U9_Z_30), .CK(clock), .Q(ops_out[30]) );
  DFF_X2 adr_2_op_reg_25_ ( .D(U7_Z_25), .CK(clock), .Q(U6_B_25_), .QN(n641)
         );
  DFF_X2 adr_2_op_reg_26_ ( .D(U7_Z_26), .CK(clock), .Q(U6_B_26_), .QN(n1300)
         );
  DFF_X2 adr_1_op_reg_31_ ( .D(U8_Z_31), .CK(clock), .Q(U6_A_31_) );
  DFF_X2 ops_out_reg_31_ ( .D(U9_Z_31), .CK(clock), .Q(ops_out[31]) );
  DFF_X2 adr_2_op_reg_31_ ( .D(U7_Z_31), .CK(clock), .Q(U6_B_31_) );
  NOR2_X4 U170 ( .A1(net4704), .A2(n759), .ZN(n695) );
  INV_X2 U171 ( .A(n878), .ZN(n648) );
  INV_X4 U172 ( .A(n846), .ZN(n1127) );
  NOR2_X4 U173 ( .A1(n846), .A2(n1129), .ZN(n840) );
  INV_X2 U174 ( .A(n647), .ZN(n777) );
  INV_X2 U175 ( .A(n785), .ZN(n786) );
  NOR2_X2 U176 ( .A1(n1260), .A2(n1261), .ZN(net4954) );
  NOR2_X2 U177 ( .A1(n831), .A2(n1183), .ZN(n842) );
  OR2_X4 U178 ( .A1(in2[0]), .A2(in4[29]), .ZN(n758) );
  AND2_X4 U179 ( .A1(n741), .A2(n717), .ZN(n630) );
  NAND2_X2 U180 ( .A1(n624), .A2(n625), .ZN(n690) );
  NAND2_X2 U181 ( .A1(n626), .A2(n627), .ZN(n680) );
  NAND2_X2 U182 ( .A1(n628), .A2(n629), .ZN(n670) );
  NAND2_X2 U183 ( .A1(n1044), .A2(in4[4]), .ZN(n1045) );
  OAI21_X2 U184 ( .B1(n891), .B2(in2[4]), .A(n812), .ZN(n997) );
  XNOR2_X1 U185 ( .A(n985), .B(in4[0]), .ZN(n980) );
  AND3_X4 U186 ( .A1(net3546), .A2(n753), .A3(n659), .ZN(n769) );
  NOR2_X2 U187 ( .A1(n1181), .A2(n1182), .ZN(n843) );
  OAI22_X2 U188 ( .A1(n905), .A2(n884), .B1(n1191), .B2(n883), .ZN(n666) );
  OAI22_X2 U189 ( .A1(n717), .A2(net3677), .B1(n630), .B2(n728), .ZN(net3640)
         );
  NAND2_X2 U190 ( .A1(n631), .A2(n632), .ZN(n676) );
  NAND2_X2 U191 ( .A1(n633), .A2(n634), .ZN(n671) );
  NAND2_X2 U192 ( .A1(n635), .A2(n636), .ZN(n669) );
  NAND2_X2 U193 ( .A1(n637), .A2(n638), .ZN(n663) );
  OAI22_X2 U194 ( .A1(in4[25]), .A2(in2[28]), .B1(in4[26]), .B2(in2[29]), .ZN(
        n726) );
  OAI21_X2 U195 ( .B1(n639), .B2(in3[12]), .A(n709), .ZN(n698) );
  INV_X4 U196 ( .A(net5590), .ZN(n639) );
  NAND3_X2 U197 ( .A1(n640), .A2(n767), .A3(n1063), .ZN(n897) );
  INV_X4 U198 ( .A(in4[6]), .ZN(n640) );
  XNOR2_X2 U199 ( .A(in4[4]), .B(n1047), .ZN(n1034) );
  XNOR2_X2 U200 ( .A(in4[2]), .B(n1015), .ZN(n998) );
  NAND3_X1 U201 ( .A1(n739), .A2(n735), .A3(net5243), .ZN(n743) );
  XNOR2_X2 U202 ( .A(in1[20]), .B(in1[18]), .ZN(n982) );
  NAND2_X2 U203 ( .A1(n641), .A2(n642), .ZN(n681) );
  NAND2_X2 U204 ( .A1(n643), .A2(n644), .ZN(n675) );
  NAND2_X2 U205 ( .A1(n645), .A2(n646), .ZN(n668) );
  AOI21_X2 U206 ( .B1(n717), .B2(n741), .A(n728), .ZN(n724) );
  OAI21_X1 U207 ( .B1(n696), .B2(n1158), .A(n818), .ZN(n647) );
  NAND3_X2 U208 ( .A1(net5590), .A2(n792), .A3(n791), .ZN(n797) );
  OAI22_X2 U209 ( .A1(n773), .A2(n1105), .B1(n1107), .B2(n1106), .ZN(n774) );
  XNOR2_X2 U210 ( .A(n1048), .B(in2[8]), .ZN(n662) );
  NAND3_X1 U211 ( .A1(n890), .A2(n889), .A3(in2[3]), .ZN(n886) );
  XNOR2_X1 U212 ( .A(n1029), .B(n1016), .ZN(n1017) );
  NOR3_X2 U213 ( .A1(n842), .A2(n843), .A3(in4[17]), .ZN(n1193) );
  NAND2_X2 U214 ( .A1(n648), .A2(in4[13]), .ZN(n818) );
  OAI22_X2 U215 ( .A1(n1057), .A2(n1058), .B1(n1060), .B2(n1059), .ZN(n1070)
         );
  NAND2_X2 U216 ( .A1(n649), .A2(n650), .ZN(n674) );
  OAI211_X1 U217 ( .C1(n651), .C2(n745), .A(n718), .B(n719), .ZN(net3677) );
  INV_X4 U218 ( .A(net3683), .ZN(n651) );
  OR2_X4 U219 ( .A1(in1[28]), .A2(in3[18]), .ZN(net4701) );
  OR2_X4 U220 ( .A1(net3997), .A2(n787), .ZN(n795) );
  XOR2_X2 U221 ( .A(in1[26]), .B(in1[24]), .Z(net4826) );
  NAND3_X2 U222 ( .A1(n969), .A2(n968), .A3(in3[0]), .ZN(n778) );
  XOR2_X2 U223 ( .A(n1314), .B(n930), .Z(n1315) );
  XOR2_X2 U224 ( .A(n1302), .B(n935), .Z(n1303) );
  XOR2_X2 U225 ( .A(n1170), .B(n947), .Z(n1171) );
  XNOR2_X2 U226 ( .A(n826), .B(n861), .ZN(n1231) );
  XOR2_X1 U227 ( .A(n774), .B(n870), .Z(n1108) );
  XOR2_X1 U228 ( .A(n896), .B(n1078), .Z(n1079) );
  XNOR2_X1 U229 ( .A(n1062), .B(n1049), .ZN(n1050) );
  XNOR2_X2 U230 ( .A(in4[3]), .B(n1032), .ZN(n1016) );
  OAI21_X2 U231 ( .B1(in4[24]), .B2(n719), .A(n743), .ZN(n652) );
  INV_X4 U232 ( .A(n652), .ZN(n736) );
  NAND2_X2 U233 ( .A1(in1[7]), .A2(in3[29]), .ZN(n838) );
  NOR2_X2 U234 ( .A1(n1175), .A2(n1176), .ZN(n845) );
  NOR2_X2 U235 ( .A1(n833), .A2(n840), .ZN(n835) );
  XNOR2_X2 U236 ( .A(in1[25]), .B(in1[27]), .ZN(n1086) );
  XOR2_X2 U237 ( .A(in1[25]), .B(in1[23]), .Z(net4544) );
  XOR2_X2 U238 ( .A(n982), .B(in1[11]), .Z(n990) );
  XOR2_X2 U239 ( .A(n1285), .B(n938), .Z(n1286) );
  XOR2_X2 U240 ( .A(n1268), .B(n940), .Z(n1269) );
  XOR2_X2 U241 ( .A(n1242), .B(n942), .Z(n1243) );
  XOR2_X2 U242 ( .A(n1211), .B(n945), .Z(n1212) );
  XOR2_X2 U243 ( .A(n1189), .B(n943), .Z(n1190) );
  XOR2_X2 U244 ( .A(n1154), .B(n951), .Z(n1155) );
  OAI21_X2 U245 ( .B1(n723), .B2(n726), .A(n740), .ZN(n653) );
  INV_X4 U246 ( .A(n653), .ZN(n770) );
  XOR2_X2 U247 ( .A(n819), .B(n911), .Z(n1292) );
  AND3_X4 U248 ( .A1(n707), .A2(n705), .A3(n706), .ZN(n702) );
  XOR2_X2 U249 ( .A(n788), .B(in3[11]), .Z(net4804) );
  XNOR2_X2 U250 ( .A(in4[7]), .B(n1091), .ZN(n1078) );
  XNOR2_X2 U251 ( .A(n1044), .B(n1034), .ZN(n1035) );
  XNOR2_X2 U252 ( .A(n1012), .B(n998), .ZN(n999) );
  AOI211_X2 U253 ( .C1(net3544), .C2(net5800), .A(n1317), .B(n769), .ZN(
        U7_Z_30) );
  NOR2_X2 U254 ( .A1(n834), .A2(n841), .ZN(n1139) );
  NOR2_X2 U255 ( .A1(n832), .A2(n1128), .ZN(n841) );
  OR2_X4 U256 ( .A1(n695), .A2(net4887), .ZN(n654) );
  INV_X2 U257 ( .A(n1262), .ZN(n836) );
  AOI22_X1 U258 ( .A1(n1084), .A2(in3[7]), .B1(n965), .B2(n932), .ZN(n964) );
  AOI21_X2 U259 ( .B1(net5301), .B2(n673), .A(n665), .ZN(net4920) );
  NAND2_X2 U260 ( .A1(n836), .A2(in4[22]), .ZN(net5243) );
  NOR2_X2 U261 ( .A1(n1127), .A2(in4[10]), .ZN(n832) );
  NOR2_X2 U262 ( .A1(n1005), .A2(in3[2]), .ZN(n1006) );
  OAI21_X2 U263 ( .B1(in2[28]), .B2(in4[25]), .A(net3640), .ZN(net3639) );
  AOI22_X2 U264 ( .A1(U6_A_29_), .A2(U6_B_29_), .B1(n1314), .B2(n690), .ZN(
        n926) );
  AOI22_X2 U265 ( .A1(U6_A_23_), .A2(U6_B_23_), .B1(n1268), .B2(n680), .ZN(
        n919) );
  AOI22_X2 U266 ( .A1(U6_A_21_), .A2(U6_B_21_), .B1(n1242), .B2(n676), .ZN(
        n918) );
  AOI22_X2 U267 ( .A1(U6_A_19_), .A2(U6_B_19_), .B1(n1211), .B2(n675), .ZN(
        n917) );
  OAI21_X2 U268 ( .B1(net3677), .B2(n717), .A(net3620), .ZN(n725) );
  AOI22_X2 U269 ( .A1(in1[26]), .A2(in3[16]), .B1(net5294), .B2(n906), .ZN(
        n905) );
  OAI21_X2 U270 ( .B1(n700), .B2(n701), .A(n672), .ZN(net5301) );
  NAND3_X2 U271 ( .A1(n698), .A2(n699), .A3(net5228), .ZN(n697) );
  NOR2_X2 U272 ( .A1(n800), .A2(n976), .ZN(n801) );
  INV_X4 U273 ( .A(n758), .ZN(net5801) );
  BUF_X4 U274 ( .A(n900), .Z(n810) );
  INV_X4 U275 ( .A(n878), .ZN(n1156) );
  NOR2_X2 U276 ( .A1(n1156), .A2(in4[13]), .ZN(n696) );
  AOI22_X2 U277 ( .A1(in1[8]), .A2(in3[30]), .B1(n882), .B2(n693), .ZN(n907)
         );
  INV_X4 U278 ( .A(n811), .ZN(n1118) );
  AOI22_X2 U279 ( .A1(in1[1]), .A2(in3[23]), .B1(n1257), .B2(n679), .ZN(n904)
         );
  NOR2_X2 U280 ( .A1(n809), .A2(in3[1]), .ZN(n989) );
  AOI22_X2 U281 ( .A1(U6_A_25_), .A2(U6_B_25_), .B1(n1285), .B2(n681), .ZN(
        n920) );
  AOI22_X2 U282 ( .A1(U6_A_27_), .A2(U6_B_27_), .B1(n1302), .B2(n689), .ZN(
        n922) );
  AOI22_X2 U283 ( .A1(U6_A_15_), .A2(U6_B_15_), .B1(n1170), .B2(n671), .ZN(
        n910) );
  AOI22_X2 U284 ( .A1(U6_A_17_), .A2(U6_B_17_), .B1(n1189), .B2(n674), .ZN(
        n916) );
  NOR2_X2 U285 ( .A1(n657), .A2(n658), .ZN(n655) );
  NAND2_X2 U286 ( .A1(n818), .A2(n656), .ZN(n658) );
  INV_X4 U287 ( .A(in4[14]), .ZN(n656) );
  NOR2_X2 U288 ( .A1(n658), .A2(n657), .ZN(n1163) );
  NOR2_X2 U289 ( .A1(n1157), .A2(n1158), .ZN(n657) );
  NOR2_X4 U290 ( .A1(n695), .A2(net4887), .ZN(n659) );
  INV_X1 U291 ( .A(n768), .ZN(n660) );
  INV_X4 U292 ( .A(n660), .ZN(n661) );
  AOI22_X2 U293 ( .A1(U6_A_13_), .A2(U6_B_13_), .B1(n1154), .B2(n670), .ZN(
        n909) );
  NOR2_X2 U294 ( .A1(n775), .A2(in4[15]), .ZN(n1175) );
  INV_X1 U295 ( .A(n1135), .ZN(n1144) );
  AOI22_X2 U296 ( .A1(U6_A_11_), .A2(U6_B_11_), .B1(n1135), .B2(n668), .ZN(
        n908) );
  INV_X1 U297 ( .A(n1054), .ZN(n1068) );
  AOI22_X2 U298 ( .A1(U6_A_5_), .A2(U6_B_5_), .B1(n1054), .B2(n667), .ZN(n925)
         );
  INV_X1 U299 ( .A(n1021), .ZN(n1036) );
  AOI22_X2 U300 ( .A1(U6_A_3_), .A2(U6_B_3_), .B1(n1021), .B2(n663), .ZN(n924)
         );
  INV_X1 U301 ( .A(n1112), .ZN(n1124) );
  AOI22_X2 U302 ( .A1(U6_A_9_), .A2(U6_B_9_), .B1(n1112), .B2(n669), .ZN(n915)
         );
  INV_X4 U303 ( .A(n778), .ZN(n809) );
  INV_X1 U304 ( .A(n1257), .ZN(n1270) );
  XNOR2_X2 U305 ( .A(n1065), .B(in2[9]), .ZN(n664) );
  AND2_X4 U306 ( .A1(in1[25]), .A2(in3[15]), .ZN(n665) );
  OR2_X4 U307 ( .A1(U6_B_5_), .A2(U6_A_5_), .ZN(n667) );
  AOI22_X2 U308 ( .A1(in1[28]), .A2(in3[18]), .B1(n666), .B2(net4701), .ZN(
        n899) );
  OR2_X4 U309 ( .A1(n704), .A2(n703), .ZN(n672) );
  OR2_X4 U310 ( .A1(in3[15]), .A2(in1[25]), .ZN(n673) );
  OR2_X4 U311 ( .A1(in3[21]), .A2(in1[31]), .ZN(n677) );
  XOR2_X2 U312 ( .A(net3997), .B(in3[10]), .Z(n678) );
  OR2_X4 U313 ( .A1(in3[23]), .A2(in1[1]), .ZN(n679) );
  AND2_X4 U314 ( .A1(n726), .A2(n740), .ZN(n682) );
  OR2_X4 U315 ( .A1(in3[26]), .A2(in1[4]), .ZN(n683) );
  XNOR2_X2 U316 ( .A(in3[30]), .B(in1[8]), .ZN(n684) );
  OR2_X4 U317 ( .A1(in4[27]), .A2(in2[30]), .ZN(n685) );
  XOR2_X2 U318 ( .A(in1[28]), .B(in3[18]), .Z(n686) );
  XOR2_X2 U319 ( .A(n704), .B(n703), .Z(n687) );
  XOR2_X2 U320 ( .A(n712), .B(n710), .Z(n688) );
  OR2_X4 U321 ( .A1(U6_B_27_), .A2(U6_A_27_), .ZN(n689) );
  OR2_X4 U322 ( .A1(in3[29]), .A2(in1[7]), .ZN(n691) );
  OR2_X4 U323 ( .A1(in3[27]), .A2(in1[5]), .ZN(n692) );
  OR2_X4 U324 ( .A1(in3[30]), .A2(in1[8]), .ZN(n693) );
  NOR2_X1 U325 ( .A1(n842), .A2(n843), .ZN(n694) );
  NOR2_X2 U326 ( .A1(net4704), .A2(n759), .ZN(n760) );
  AOI22_X4 U327 ( .A1(in2[30]), .A2(in4[27]), .B1(net5325), .B2(n685), .ZN(
        net4704) );
  NOR2_X2 U328 ( .A1(n1156), .A2(in4[13]), .ZN(n1157) );
  INV_X4 U329 ( .A(in3[14]), .ZN(n703) );
  XNOR2_X2 U330 ( .A(in1[24]), .B(in1[31]), .ZN(n704) );
  XNOR2_X2 U331 ( .A(n702), .B(n687), .ZN(net3916) );
  XNOR2_X2 U332 ( .A(n688), .B(n697), .ZN(net3941) );
  NAND2_X2 U333 ( .A1(n705), .A2(n706), .ZN(n700) );
  NAND2_X2 U334 ( .A1(n707), .A2(n708), .ZN(n701) );
  INV_X4 U335 ( .A(net3947), .ZN(n709) );
  INV_X4 U336 ( .A(in3[13]), .ZN(n710) );
  NAND2_X2 U337 ( .A1(n709), .A2(net6111), .ZN(n699) );
  INV_X4 U338 ( .A(n697), .ZN(n711) );
  NAND2_X2 U339 ( .A1(n712), .A2(n710), .ZN(n706) );
  NAND2_X2 U340 ( .A1(n712), .A2(n711), .ZN(n705) );
  NAND2_X2 U341 ( .A1(n704), .A2(n703), .ZN(n708) );
  NAND2_X2 U342 ( .A1(n711), .A2(n710), .ZN(n707) );
  XNOR2_X2 U343 ( .A(in1[23]), .B(in1[30]), .ZN(n712) );
  NOR2_X1 U344 ( .A1(n973), .A2(n1309), .ZN(U8_Z_29) );
  NOR2_X2 U345 ( .A1(n730), .A2(n731), .ZN(n729) );
  NAND2_X2 U346 ( .A1(n1174), .A2(in4[15]), .ZN(n713) );
  AOI22_X2 U347 ( .A1(in1[5]), .A2(in3[27]), .B1(n823), .B2(n692), .ZN(n902)
         );
  NAND2_X2 U348 ( .A1(n713), .A2(n1183), .ZN(n830) );
  INV_X1 U349 ( .A(n994), .ZN(n714) );
  INV_X4 U350 ( .A(n714), .ZN(n715) );
  INV_X4 U351 ( .A(n993), .ZN(n994) );
  NAND3_X1 U352 ( .A1(n718), .A2(n719), .A3(n742), .ZN(n741) );
  INV_X4 U353 ( .A(n902), .ZN(n803) );
  INV_X2 U354 ( .A(n804), .ZN(n1009) );
  INV_X1 U355 ( .A(n1070), .ZN(n1074) );
  INV_X1 U356 ( .A(n666), .ZN(n716) );
  INV_X1 U357 ( .A(n797), .ZN(net3945) );
  AND2_X2 U358 ( .A1(n907), .A2(n851), .ZN(n807) );
  NAND2_X2 U359 ( .A1(n791), .A2(n792), .ZN(net6111) );
  INV_X4 U360 ( .A(net5243), .ZN(net5018) );
  INV_X1 U361 ( .A(n790), .ZN(net5277) );
  AOI21_X4 U362 ( .B1(n720), .B2(n721), .A(n682), .ZN(net5325) );
  INV_X4 U363 ( .A(in4[24]), .ZN(n717) );
  INV_X4 U364 ( .A(net3620), .ZN(n722) );
  NOR2_X2 U365 ( .A1(n724), .A2(n725), .ZN(n723) );
  INV_X4 U366 ( .A(in4[26]), .ZN(n727) );
  NAND2_X2 U367 ( .A1(net3683), .A2(n732), .ZN(n719) );
  XNOR2_X2 U368 ( .A(in2[27]), .B(in2[31]), .ZN(n728) );
  XNOR2_X2 U369 ( .A(n728), .B(n717), .ZN(net4626) );
  XNOR2_X2 U370 ( .A(in2[16]), .B(in2[27]), .ZN(net4035) );
  XNOR2_X2 U371 ( .A(in2[17]), .B(in2[28]), .ZN(net4010) );
  XNOR2_X2 U372 ( .A(in2[29]), .B(n727), .ZN(net3637) );
  NAND2_X2 U373 ( .A1(n718), .A2(n719), .ZN(n730) );
  NAND2_X2 U374 ( .A1(n734), .A2(in4[24]), .ZN(n731) );
  NOR2_X2 U375 ( .A1(in4[24]), .A2(in4[23]), .ZN(n735) );
  NOR2_X2 U376 ( .A1(n738), .A2(n728), .ZN(n737) );
  NOR2_X2 U377 ( .A1(n722), .A2(net4724), .ZN(n721) );
  INV_X4 U378 ( .A(in4[23]), .ZN(n732) );
  NAND2_X2 U379 ( .A1(in2[29]), .A2(in4[26]), .ZN(n740) );
  INV_X4 U380 ( .A(n740), .ZN(net4724) );
  NAND2_X2 U381 ( .A1(n733), .A2(net5243), .ZN(n718) );
  NAND2_X2 U382 ( .A1(net3683), .A2(n746), .ZN(n742) );
  NAND2_X2 U383 ( .A1(net5011), .A2(net3683), .ZN(n734) );
  NAND3_X2 U384 ( .A1(net3683), .A2(net5011), .A3(n717), .ZN(n744) );
  INV_X4 U385 ( .A(n744), .ZN(n738) );
  INV_X4 U386 ( .A(n745), .ZN(n746) );
  INV_X1 U387 ( .A(net5011), .ZN(n745) );
  AOI21_X2 U388 ( .B1(n737), .B2(n736), .A(n729), .ZN(n720) );
  INV_X1 U389 ( .A(net4954), .ZN(n739) );
  NOR2_X1 U390 ( .A1(net4954), .A2(in4[23]), .ZN(n733) );
  OAI33_X1 U391 ( .A1(n761), .A2(n748), .A3(n749), .B1(n763), .B2(n750), .B3(
        n751), .ZN(n747) );
  NOR2_X2 U392 ( .A1(n747), .A2(net3512), .ZN(U7_Z_31) );
  INV_X4 U393 ( .A(n752), .ZN(n750) );
  NAND2_X2 U394 ( .A1(n764), .A2(n765), .ZN(n763) );
  OR2_X1 U395 ( .A1(net3549), .A2(n758), .ZN(n765) );
  OR2_X1 U396 ( .A1(net4887), .A2(net3549), .ZN(n766) );
  OR2_X4 U397 ( .A1(n760), .A2(n766), .ZN(n764) );
  INV_X4 U398 ( .A(n751), .ZN(n749) );
  NOR2_X2 U399 ( .A1(n749), .A2(n752), .ZN(n754) );
  OAI22_X2 U400 ( .A1(n749), .A2(net3525), .B1(n748), .B2(n754), .ZN(net3523)
         );
  INV_X4 U401 ( .A(net3525), .ZN(n748) );
  NAND2_X2 U402 ( .A1(n762), .A2(n753), .ZN(n761) );
  INV_X4 U403 ( .A(net5800), .ZN(n762) );
  XNOR2_X2 U404 ( .A(in4[31]), .B(in2[2]), .ZN(n751) );
  NAND2_X2 U405 ( .A1(n755), .A2(n756), .ZN(n752) );
  INV_X4 U406 ( .A(in4[30]), .ZN(n756) );
  INV_X4 U407 ( .A(in2[1]), .ZN(n755) );
  XOR2_X2 U408 ( .A(n755), .B(in4[30]), .Z(net3546) );
  NOR2_X2 U409 ( .A1(net3544), .A2(n758), .ZN(n757) );
  NAND2_X2 U410 ( .A1(in4[29]), .A2(in2[0]), .ZN(n753) );
  INV_X4 U411 ( .A(n753), .ZN(net3549) );
  OAI22_X2 U412 ( .A1(net3544), .A2(n753), .B1(net3549), .B2(n757), .ZN(
        net3548) );
  NOR2_X2 U413 ( .A1(in4[28]), .A2(in2[31]), .ZN(n759) );
  NOR2_X1 U414 ( .A1(n832), .A2(n1128), .ZN(n833) );
  XOR2_X2 U415 ( .A(n654), .B(n895), .Z(n1310) );
  NOR2_X2 U416 ( .A1(n659), .A2(net5801), .ZN(net5800) );
  INV_X1 U417 ( .A(net3999), .ZN(net5364) );
  NAND2_X2 U418 ( .A1(n780), .A2(n662), .ZN(n767) );
  NAND2_X2 U419 ( .A1(n780), .A2(n662), .ZN(n781) );
  NAND2_X2 U420 ( .A1(n781), .A2(n1063), .ZN(n768) );
  INV_X1 U421 ( .A(net3546), .ZN(net3544) );
  INV_X4 U422 ( .A(n985), .ZN(n776) );
  NAND2_X2 U423 ( .A1(n797), .A2(in3[12]), .ZN(net5228) );
  AND2_X4 U424 ( .A1(n768), .A2(in4[6]), .ZN(n898) );
  NAND2_X2 U425 ( .A1(n801), .A2(n972), .ZN(n969) );
  INV_X4 U426 ( .A(n1064), .ZN(n780) );
  INV_X1 U427 ( .A(n1174), .ZN(n771) );
  INV_X1 U428 ( .A(n1098), .ZN(n772) );
  NOR2_X1 U429 ( .A1(n1103), .A2(in4[8]), .ZN(n773) );
  NOR2_X2 U430 ( .A1(n1103), .A2(in4[8]), .ZN(n1104) );
  OAI22_X2 U431 ( .A1(n777), .A2(n656), .B1(n1163), .B2(n1164), .ZN(n775) );
  NOR2_X2 U432 ( .A1(n1070), .A2(in3[6]), .ZN(n1071) );
  NAND2_X1 U433 ( .A1(n779), .A2(n776), .ZN(n995) );
  AND2_X4 U434 ( .A1(in4[0]), .A2(in4[1]), .ZN(n779) );
  NOR2_X4 U435 ( .A1(n1062), .A2(in4[5]), .ZN(n1064) );
  NAND2_X1 U436 ( .A1(n1062), .A2(in4[5]), .ZN(n1063) );
  NOR2_X4 U437 ( .A1(n994), .A2(in4[1]), .ZN(n996) );
  NAND2_X1 U438 ( .A1(in2[19]), .A2(n822), .ZN(n783) );
  NAND2_X2 U439 ( .A1(n782), .A2(in2[8]), .ZN(n784) );
  NAND2_X2 U440 ( .A1(n783), .A2(n784), .ZN(n891) );
  INV_X2 U441 ( .A(in2[19]), .ZN(n782) );
  INV_X2 U442 ( .A(in2[8]), .ZN(n822) );
  NAND2_X2 U443 ( .A1(n891), .A2(in2[4]), .ZN(n812) );
  INV_X2 U444 ( .A(n1103), .ZN(n1107) );
  INV_X1 U445 ( .A(n694), .ZN(n785) );
  NOR2_X2 U446 ( .A1(n1114), .A2(in3[9]), .ZN(n1115) );
  NOR2_X2 U447 ( .A1(n1038), .A2(in3[4]), .ZN(n1039) );
  NOR2_X4 U448 ( .A1(n1044), .A2(in4[4]), .ZN(n1046) );
  INV_X4 U449 ( .A(in3[10]), .ZN(n787) );
  XNOR2_X2 U450 ( .A(n789), .B(net5579), .ZN(n788) );
  XNOR2_X2 U451 ( .A(in1[21]), .B(in1[23]), .ZN(net4627) );
  XNOR2_X2 U452 ( .A(in1[21]), .B(net4311), .ZN(net4221) );
  XNOR2_X2 U453 ( .A(in1[28]), .B(in1[26]), .ZN(net4044) );
  NAND2_X2 U454 ( .A1(in3[11]), .A2(n790), .ZN(net5590) );
  INV_X4 U455 ( .A(in1[30]), .ZN(net5579) );
  NAND2_X2 U456 ( .A1(net3997), .A2(n787), .ZN(n793) );
  NAND2_X2 U457 ( .A1(net3999), .A2(n793), .ZN(n794) );
  NAND2_X2 U458 ( .A1(n794), .A2(n795), .ZN(n790) );
  NAND2_X2 U459 ( .A1(n790), .A2(n796), .ZN(n792) );
  NAND2_X2 U460 ( .A1(n796), .A2(in3[11]), .ZN(n791) );
  INV_X4 U461 ( .A(n788), .ZN(n796) );
  XNOR2_X2 U462 ( .A(in1[28]), .B(in1[21]), .ZN(n789) );
  INV_X1 U463 ( .A(n1288), .ZN(n798) );
  INV_X1 U464 ( .A(n798), .ZN(n799) );
  NAND2_X2 U465 ( .A1(n979), .A2(n978), .ZN(n885) );
  NOR2_X2 U466 ( .A1(n1098), .A2(in3[8]), .ZN(n1099) );
  INV_X2 U467 ( .A(n971), .ZN(n800) );
  NAND2_X2 U468 ( .A1(n972), .A2(n971), .ZN(n802) );
  NAND2_X2 U469 ( .A1(in1[17]), .A2(in1[19]), .ZN(n971) );
  OAI22_X1 U470 ( .A1(n778), .A2(n991), .B1(n990), .B2(n989), .ZN(n804) );
  INV_X1 U471 ( .A(in1[18]), .ZN(n805) );
  NAND2_X1 U472 ( .A1(n691), .A2(n827), .ZN(n806) );
  XNOR2_X2 U473 ( .A(n903), .B(n684), .ZN(n1316) );
  NOR2_X2 U474 ( .A1(n807), .A2(n808), .ZN(U8_Z_31) );
  NAND2_X2 U475 ( .A1(n817), .A2(n975), .ZN(n808) );
  OR2_X4 U476 ( .A1(n1146), .A2(in4[12]), .ZN(n881) );
  INV_X2 U477 ( .A(n1056), .ZN(n1060) );
  INV_X1 U478 ( .A(in3[5]), .ZN(n1059) );
  NOR2_X2 U479 ( .A1(n1029), .A2(in4[3]), .ZN(n1031) );
  OR2_X2 U480 ( .A1(n840), .A2(in4[11]), .ZN(n834) );
  OAI22_X1 U481 ( .A1(n772), .A2(n1101), .B1(n1099), .B2(n1100), .ZN(n811) );
  INV_X4 U482 ( .A(net4920), .ZN(net5294) );
  INV_X4 U483 ( .A(n901), .ZN(n823) );
  NAND2_X2 U484 ( .A1(n806), .A2(n838), .ZN(n813) );
  NAND2_X2 U485 ( .A1(n839), .A2(n838), .ZN(n882) );
  INV_X2 U486 ( .A(n813), .ZN(n903) );
  INV_X4 U487 ( .A(n828), .ZN(n814) );
  NAND2_X2 U488 ( .A1(n815), .A2(n816), .ZN(n817) );
  INV_X4 U489 ( .A(n907), .ZN(n815) );
  INV_X4 U490 ( .A(n851), .ZN(n816) );
  INV_X1 U491 ( .A(net4704), .ZN(net5264) );
  INV_X2 U492 ( .A(net5264), .ZN(net5265) );
  XNOR2_X2 U493 ( .A(n934), .B(in2[16]), .ZN(n1158) );
  OR2_X4 U494 ( .A1(n1121), .A2(in4[9]), .ZN(n848) );
  OAI22_X1 U495 ( .A1(n1290), .A2(n1289), .B1(n1287), .B2(n799), .ZN(n819) );
  INV_X4 U496 ( .A(n849), .ZN(n827) );
  INV_X1 U497 ( .A(n1023), .ZN(n1027) );
  NAND2_X1 U498 ( .A1(in2[18]), .A2(in2[7]), .ZN(n889) );
  INV_X1 U499 ( .A(n716), .ZN(n820) );
  NOR2_X2 U500 ( .A1(n825), .A2(n845), .ZN(n831) );
  INV_X2 U501 ( .A(n1259), .ZN(n1262) );
  AOI22_X2 U502 ( .A1(in1[31]), .A2(in3[21]), .B1(n1230), .B2(n677), .ZN(n900)
         );
  AOI22_X2 U503 ( .A1(in1[6]), .A2(in3[28]), .B1(n803), .B2(n850), .ZN(n849)
         );
  XOR2_X1 U504 ( .A(n1119), .B(in1[20]), .Z(net3997) );
  INV_X4 U505 ( .A(n964), .ZN(n1098) );
  OR2_X2 U506 ( .A1(n1084), .A2(in3[7]), .ZN(n965) );
  NAND2_X2 U507 ( .A1(n802), .A2(n976), .ZN(n968) );
  NOR2_X2 U508 ( .A1(net5018), .A2(net4954), .ZN(net5011) );
  INV_X1 U509 ( .A(n887), .ZN(n821) );
  NAND2_X2 U510 ( .A1(n827), .A2(n691), .ZN(n839) );
  XOR2_X1 U511 ( .A(n997), .B(in4[1]), .Z(n986) );
  NOR2_X2 U512 ( .A1(n1012), .A2(in4[2]), .ZN(n1014) );
  INV_X1 U513 ( .A(n823), .ZN(n824) );
  AOI22_X2 U514 ( .A1(in1[4]), .A2(in3[26]), .B1(n1291), .B2(n683), .ZN(n901)
         );
  INV_X1 U515 ( .A(in2[18]), .ZN(n1165) );
  INV_X2 U516 ( .A(n713), .ZN(n825) );
  OAI21_X4 U517 ( .B1(n1046), .B2(n1047), .A(n1045), .ZN(n1062) );
  OAI22_X1 U518 ( .A1(net5579), .A2(n1229), .B1(n814), .B2(n1227), .ZN(n826)
         );
  OAI22_X2 U519 ( .A1(net5579), .A2(n1229), .B1(n1228), .B2(n1227), .ZN(n1230)
         );
  NAND2_X2 U520 ( .A1(n776), .A2(in4[0]), .ZN(n993) );
  INV_X1 U521 ( .A(n1228), .ZN(n828) );
  NOR2_X2 U522 ( .A1(n1259), .A2(in4[22]), .ZN(n1260) );
  NOR2_X4 U523 ( .A1(n829), .A2(in4[7]), .ZN(n1090) );
  INV_X4 U524 ( .A(n896), .ZN(n1088) );
  INV_X4 U525 ( .A(n896), .ZN(n829) );
  AOI21_X4 U526 ( .B1(n897), .B2(n664), .A(n898), .ZN(n896) );
  XOR2_X1 U527 ( .A(n878), .B(n1149), .Z(n1150) );
  INV_X1 U528 ( .A(n1146), .ZN(n1148) );
  INV_X1 U529 ( .A(n836), .ZN(n837) );
  OAI21_X4 U530 ( .B1(n996), .B2(n997), .A(n995), .ZN(n1012) );
  XOR2_X1 U531 ( .A(n986), .B(n715), .Z(n987) );
  OAI21_X4 U532 ( .B1(n1031), .B2(n1032), .A(n1030), .ZN(n1044) );
  NAND2_X2 U533 ( .A1(n1029), .A2(in4[3]), .ZN(n1030) );
  OAI21_X4 U534 ( .B1(n1090), .B2(n1091), .A(n1089), .ZN(n1103) );
  OAI21_X4 U535 ( .B1(n1014), .B2(n1015), .A(n1013), .ZN(n1029) );
  NAND2_X2 U536 ( .A1(n1012), .A2(in4[2]), .ZN(n1013) );
  INV_X2 U537 ( .A(in4[10]), .ZN(n1129) );
  INV_X1 U538 ( .A(in4[16]), .ZN(n1183) );
  INV_X4 U539 ( .A(n1122), .ZN(n847) );
  INV_X1 U540 ( .A(net5301), .ZN(net3875) );
  XNOR2_X1 U541 ( .A(n746), .B(n854), .ZN(n1264) );
  INV_X1 U542 ( .A(n803), .ZN(n844) );
  AOI22_X4 U543 ( .A1(n774), .A2(in4[9]), .B1(n848), .B2(n847), .ZN(n846) );
  OR2_X1 U544 ( .A1(in3[16]), .A2(in1[26]), .ZN(n906) );
  XOR2_X2 U545 ( .A(net4826), .B(in1[17]), .Z(n932) );
  XNOR2_X2 U546 ( .A(net3677), .B(net4626), .ZN(n1273) );
  INV_X4 U547 ( .A(n852), .ZN(n923) );
  INV_X4 U548 ( .A(n853), .ZN(n927) );
  INV_X4 U549 ( .A(n856), .ZN(n921) );
  OAI22_X2 U550 ( .A1(n1096), .A2(n1095), .B1(n923), .B2(n1094), .ZN(n856) );
  NOR2_X2 U551 ( .A1(net3572), .A2(net3573), .ZN(net4887) );
  NOR2_X2 U552 ( .A1(in3[17]), .A2(in1[27]), .ZN(n884) );
  XNOR2_X1 U553 ( .A(n820), .B(n686), .ZN(n1192) );
  OR2_X4 U554 ( .A1(in3[28]), .A2(in1[6]), .ZN(n850) );
  XNOR2_X1 U555 ( .A(n1184), .B(in2[9]), .ZN(n894) );
  XNOR2_X2 U556 ( .A(in3[31]), .B(in1[9]), .ZN(n851) );
  XNOR2_X1 U557 ( .A(in1[22]), .B(in1[24]), .ZN(n912) );
  XNOR2_X1 U558 ( .A(n1196), .B(in2[10]), .ZN(n892) );
  XNOR2_X1 U559 ( .A(net5265), .B(n913), .ZN(n1306) );
  XNOR2_X1 U560 ( .A(net3640), .B(n1280), .ZN(n1281) );
  XOR2_X1 U561 ( .A(in4[25]), .B(in2[28]), .Z(n1280) );
  OAI22_X2 U562 ( .A1(n1082), .A2(n1081), .B1(n925), .B2(n1080), .ZN(n852) );
  OAI22_X2 U563 ( .A1(n1003), .A2(n1002), .B1(n1001), .B2(n1000), .ZN(n853) );
  XOR2_X2 U564 ( .A(in4[23]), .B(net3683), .Z(n854) );
  XNOR2_X1 U565 ( .A(n837), .B(n855), .ZN(n1252) );
  XOR2_X2 U566 ( .A(in4[22]), .B(n1261), .Z(n855) );
  XNOR2_X1 U567 ( .A(n922), .B(n931), .ZN(n1307) );
  XNOR2_X1 U568 ( .A(n1250), .B(n857), .ZN(n1238) );
  XOR2_X2 U569 ( .A(in4[21]), .B(n1248), .Z(n857) );
  XNOR2_X1 U570 ( .A(n1223), .B(n858), .ZN(n1207) );
  XOR2_X2 U571 ( .A(in4[19]), .B(n1221), .Z(n858) );
  XNOR2_X1 U572 ( .A(n1205), .B(n859), .ZN(n1197) );
  XOR2_X2 U573 ( .A(in4[18]), .B(n1203), .Z(n859) );
  XNOR2_X1 U574 ( .A(n1236), .B(n860), .ZN(n1225) );
  XOR2_X2 U575 ( .A(in4[20]), .B(n1234), .Z(n860) );
  XNOR2_X1 U576 ( .A(n933), .B(in2[15]), .ZN(n1147) );
  XNOR2_X1 U577 ( .A(n782), .B(in2[30]), .ZN(n933) );
  XNOR2_X1 U578 ( .A(n919), .B(n937), .ZN(n1274) );
  XNOR2_X1 U579 ( .A(n920), .B(n936), .ZN(n1295) );
  XOR2_X1 U580 ( .A(in3[21]), .B(in1[31]), .Z(n861) );
  XNOR2_X1 U581 ( .A(n1184), .B(in2[31]), .ZN(n934) );
  XNOR2_X1 U582 ( .A(n831), .B(n862), .ZN(n1177) );
  XOR2_X2 U583 ( .A(in4[16]), .B(n1182), .Z(n862) );
  XNOR2_X1 U584 ( .A(n786), .B(n863), .ZN(n1185) );
  XOR2_X2 U585 ( .A(in4[17]), .B(n1194), .Z(n863) );
  XOR2_X1 U586 ( .A(in3[16]), .B(in1[26]), .Z(n1172) );
  XOR2_X1 U587 ( .A(in3[17]), .B(in1[27]), .Z(n1179) );
  XNOR2_X1 U588 ( .A(n777), .B(n864), .ZN(n1159) );
  XOR2_X2 U589 ( .A(in4[14]), .B(n1164), .Z(n864) );
  XNOR2_X1 U590 ( .A(n771), .B(n865), .ZN(n1166) );
  XOR2_X2 U591 ( .A(in4[15]), .B(n1176), .Z(n865) );
  XNOR2_X1 U592 ( .A(net5364), .B(n678), .ZN(n1120) );
  XNOR2_X1 U593 ( .A(net5277), .B(net4804), .ZN(n1126) );
  XNOR2_X1 U594 ( .A(net3945), .B(n866), .ZN(n1138) );
  XOR2_X1 U595 ( .A(in3[12]), .B(net3947), .Z(n866) );
  XNOR2_X1 U596 ( .A(n835), .B(n867), .ZN(n1131) );
  XOR2_X1 U597 ( .A(in4[11]), .B(n1140), .Z(n867) );
  XNOR2_X1 U598 ( .A(n1118), .B(n868), .ZN(n1102) );
  XOR2_X1 U599 ( .A(in3[9]), .B(n1116), .Z(n868) );
  XNOR2_X1 U600 ( .A(n1107), .B(n869), .ZN(n1093) );
  XOR2_X1 U601 ( .A(in4[8]), .B(n1105), .Z(n869) );
  XOR2_X1 U602 ( .A(in4[9]), .B(n1122), .Z(n870) );
  XNOR2_X1 U603 ( .A(n846), .B(n871), .ZN(n1123) );
  XOR2_X1 U604 ( .A(in4[10]), .B(n1128), .Z(n871) );
  XNOR2_X1 U605 ( .A(n772), .B(n872), .ZN(n1087) );
  XOR2_X1 U606 ( .A(in3[8]), .B(n1100), .Z(n872) );
  XNOR2_X1 U607 ( .A(n1074), .B(n873), .ZN(n1061) );
  XOR2_X1 U608 ( .A(in3[6]), .B(n1072), .Z(n873) );
  XNOR2_X1 U609 ( .A(n923), .B(n955), .ZN(n1083) );
  XNOR2_X1 U610 ( .A(n921), .B(n956), .ZN(n1097) );
  XNOR2_X1 U611 ( .A(n1042), .B(n874), .ZN(n1028) );
  XOR2_X1 U612 ( .A(in3[4]), .B(n1040), .Z(n874) );
  XNOR2_X1 U613 ( .A(n1060), .B(n875), .ZN(n1043) );
  XOR2_X1 U614 ( .A(in3[5]), .B(n1058), .Z(n875) );
  XOR2_X1 U615 ( .A(in4[5]), .B(n662), .Z(n1049) );
  XNOR2_X1 U616 ( .A(n661), .B(n1066), .ZN(n1067) );
  XOR2_X1 U617 ( .A(in4[6]), .B(n664), .Z(n1066) );
  XNOR2_X1 U618 ( .A(U6_B_5_), .B(U6_A_5_), .ZN(n959) );
  XNOR2_X1 U619 ( .A(n1068), .B(n959), .ZN(n1055) );
  XNOR2_X1 U620 ( .A(n1027), .B(n876), .ZN(n1011) );
  XOR2_X1 U621 ( .A(in3[3]), .B(n1025), .Z(n876) );
  XNOR2_X1 U622 ( .A(n990), .B(in3[1]), .ZN(n960) );
  XOR2_X1 U623 ( .A(n960), .B(n778), .Z(n984) );
  XNOR2_X1 U624 ( .A(U6_B_4_), .B(U6_A_4_), .ZN(n958) );
  XNOR2_X1 U625 ( .A(n924), .B(n958), .ZN(n1037) );
  XNOR2_X1 U626 ( .A(U6_B_3_), .B(U6_A_3_), .ZN(n957) );
  XNOR2_X1 U627 ( .A(n1036), .B(n957), .ZN(n1022) );
  XNOR2_X1 U628 ( .A(n1009), .B(n877), .ZN(n992) );
  XOR2_X1 U629 ( .A(in3[2]), .B(n1007), .Z(n877) );
  XOR2_X1 U630 ( .A(n983), .B(in3[0]), .Z(n977) );
  INV_X4 U631 ( .A(n1148), .ZN(n879) );
  INV_X4 U632 ( .A(n1147), .ZN(n880) );
  INV_X1 U633 ( .A(in1[27]), .ZN(n1191) );
  INV_X4 U634 ( .A(in3[17]), .ZN(n883) );
  AOI22_X4 U635 ( .A1(n879), .A2(in4[12]), .B1(n881), .B2(n880), .ZN(n878) );
  NAND2_X2 U636 ( .A1(n886), .A2(n885), .ZN(n985) );
  NAND2_X2 U637 ( .A1(n888), .A2(n887), .ZN(n890) );
  NAND2_X2 U638 ( .A1(n890), .A2(n889), .ZN(n979) );
  INV_X2 U639 ( .A(in2[7]), .ZN(n887) );
  INV_X2 U640 ( .A(in2[18]), .ZN(n888) );
  INV_X4 U641 ( .A(n975), .ZN(n973) );
  INV_X4 U642 ( .A(n975), .ZN(n974) );
  XNOR2_X2 U643 ( .A(n892), .B(in2[6]), .ZN(n1032) );
  XNOR2_X2 U644 ( .A(n893), .B(in1[13]), .ZN(n1025) );
  XNOR2_X2 U645 ( .A(n1010), .B(in1[22]), .ZN(n893) );
  XNOR2_X2 U646 ( .A(n894), .B(in2[5]), .ZN(n1015) );
  XNOR2_X2 U647 ( .A(in4[29]), .B(in2[0]), .ZN(n895) );
  XNOR2_X2 U648 ( .A(in3[26]), .B(in1[4]), .ZN(n911) );
  XOR2_X2 U649 ( .A(n912), .B(in1[15]), .Z(n1058) );
  XOR2_X2 U650 ( .A(net4627), .B(in1[14]), .Z(n1040) );
  XNOR2_X2 U651 ( .A(in4[28]), .B(in2[31]), .ZN(n913) );
  XNOR2_X2 U652 ( .A(n770), .B(n914), .ZN(n1298) );
  XNOR2_X2 U653 ( .A(in4[27]), .B(in2[30]), .ZN(n914) );
  XNOR2_X2 U654 ( .A(n799), .B(n928), .ZN(n1279) );
  XNOR2_X2 U655 ( .A(in3[25]), .B(in1[3]), .ZN(n928) );
  XNOR2_X2 U656 ( .A(n1270), .B(n929), .ZN(n1258) );
  XNOR2_X2 U657 ( .A(in3[23]), .B(in1[1]), .ZN(n929) );
  XNOR2_X2 U658 ( .A(n1086), .B(n805), .ZN(n1100) );
  XNOR2_X2 U659 ( .A(net4544), .B(in1[16]), .ZN(n1072) );
  XNOR2_X2 U660 ( .A(n966), .B(n1271), .ZN(n1272) );
  XNOR2_X2 U661 ( .A(U6_B_29_), .B(U6_A_29_), .ZN(n930) );
  XNOR2_X2 U662 ( .A(U6_B_28_), .B(U6_A_28_), .ZN(n931) );
  XNOR2_X2 U663 ( .A(U6_B_27_), .B(U6_A_27_), .ZN(n935) );
  XNOR2_X2 U664 ( .A(U6_B_26_), .B(U6_A_26_), .ZN(n936) );
  XNOR2_X2 U665 ( .A(U6_B_24_), .B(U6_A_24_), .ZN(n937) );
  XNOR2_X2 U666 ( .A(U6_B_25_), .B(U6_A_25_), .ZN(n938) );
  XNOR2_X2 U667 ( .A(n918), .B(n939), .ZN(n1253) );
  XNOR2_X2 U668 ( .A(U6_B_22_), .B(U6_A_22_), .ZN(n939) );
  XNOR2_X2 U669 ( .A(U6_B_23_), .B(U6_A_23_), .ZN(n940) );
  XNOR2_X2 U670 ( .A(net4304), .B(n1172), .ZN(n1173) );
  XNOR2_X2 U671 ( .A(n967), .B(n1179), .ZN(n1180) );
  XNOR2_X2 U672 ( .A(n917), .B(n941), .ZN(n1226) );
  XNOR2_X2 U673 ( .A(U6_B_20_), .B(U6_A_20_), .ZN(n941) );
  XNOR2_X2 U674 ( .A(U6_B_21_), .B(U6_A_21_), .ZN(n942) );
  XNOR2_X2 U675 ( .A(U6_B_17_), .B(U6_A_17_), .ZN(n943) );
  XNOR2_X2 U676 ( .A(n916), .B(n944), .ZN(n1198) );
  XNOR2_X2 U677 ( .A(U6_B_18_), .B(U6_A_18_), .ZN(n944) );
  XNOR2_X2 U678 ( .A(U6_B_19_), .B(U6_A_19_), .ZN(n945) );
  XNOR2_X2 U679 ( .A(in4[12]), .B(n1147), .ZN(n1142) );
  XNOR2_X2 U680 ( .A(n909), .B(n946), .ZN(n1160) );
  XNOR2_X2 U681 ( .A(U6_B_14_), .B(U6_A_14_), .ZN(n946) );
  XNOR2_X2 U682 ( .A(U6_B_15_), .B(U6_A_15_), .ZN(n947) );
  XNOR2_X2 U683 ( .A(n910), .B(n948), .ZN(n1178) );
  XNOR2_X2 U684 ( .A(U6_B_16_), .B(U6_A_16_), .ZN(n948) );
  XNOR2_X2 U685 ( .A(in4[13]), .B(n1158), .ZN(n1149) );
  XNOR2_X2 U686 ( .A(n1144), .B(n949), .ZN(n1136) );
  XNOR2_X2 U687 ( .A(U6_B_11_), .B(U6_A_11_), .ZN(n949) );
  XNOR2_X2 U688 ( .A(n908), .B(n950), .ZN(n1145) );
  XNOR2_X2 U689 ( .A(U6_B_12_), .B(U6_A_12_), .ZN(n950) );
  XNOR2_X2 U690 ( .A(U6_B_13_), .B(U6_A_13_), .ZN(n951) );
  XNOR2_X2 U691 ( .A(n1124), .B(n952), .ZN(n1113) );
  XNOR2_X2 U692 ( .A(U6_B_9_), .B(U6_A_9_), .ZN(n952) );
  XNOR2_X2 U693 ( .A(n915), .B(n953), .ZN(n1125) );
  XNOR2_X2 U694 ( .A(U6_B_10_), .B(U6_A_10_), .ZN(n953) );
  XNOR2_X2 U695 ( .A(n925), .B(n954), .ZN(n1069) );
  XNOR2_X2 U696 ( .A(U6_B_6_), .B(U6_A_6_), .ZN(n954) );
  XNOR2_X2 U697 ( .A(U6_B_7_), .B(U6_A_7_), .ZN(n955) );
  XNOR2_X2 U698 ( .A(U6_B_8_), .B(U6_A_8_), .ZN(n956) );
  AND2_X1 U699 ( .A1(n980), .A2(n975), .ZN(n961) );
  XNOR2_X2 U700 ( .A(n927), .B(n962), .ZN(n1004) );
  XNOR2_X2 U701 ( .A(U6_B_2_), .B(U6_A_2_), .ZN(n962) );
  XOR2_X2 U702 ( .A(n963), .B(n1000), .Z(n988) );
  XOR2_X2 U703 ( .A(U6_B_1_), .B(U6_A_1_), .Z(n963) );
  INV_X4 U704 ( .A(reset), .ZN(n975) );
  XOR2_X1 U705 ( .A(n810), .B(n1244), .Z(n1245) );
  XOR2_X1 U706 ( .A(n1085), .B(n1075), .Z(n1076) );
  INV_X1 U707 ( .A(n1084), .ZN(n1085) );
  INV_X1 U708 ( .A(n1038), .ZN(n1042) );
  INV_X1 U709 ( .A(n1201), .ZN(n1205) );
  NOR2_X2 U710 ( .A1(n1023), .A2(in3[3]), .ZN(n1024) );
  INV_X1 U711 ( .A(n1219), .ZN(n1223) );
  INV_X1 U712 ( .A(n1232), .ZN(n1236) );
  INV_X1 U713 ( .A(n1246), .ZN(n1250) );
  INV_X1 U714 ( .A(n904), .ZN(n966) );
  INV_X1 U715 ( .A(net4311), .ZN(net4335) );
  INV_X2 U716 ( .A(in1[19]), .ZN(net4311) );
  INV_X1 U717 ( .A(n905), .ZN(n967) );
  INV_X1 U718 ( .A(in1[20]), .ZN(n1010) );
  INV_X1 U719 ( .A(net4920), .ZN(net4304) );
  NAND2_X2 U720 ( .A1(n969), .A2(n968), .ZN(n983) );
  NAND2_X2 U721 ( .A1(n970), .A2(net4311), .ZN(n972) );
  INV_X2 U722 ( .A(in1[17]), .ZN(n970) );
  XOR2_X1 U723 ( .A(n824), .B(n1296), .Z(n1297) );
  XOR2_X1 U724 ( .A(n844), .B(n1304), .Z(n1305) );
  XOR2_X1 U725 ( .A(n849), .B(n1308), .Z(n1309) );
  XOR2_X1 U726 ( .A(net3875), .B(n1161), .Z(n1162) );
  XOR2_X1 U727 ( .A(n899), .B(n1199), .Z(n1200) );
  XOR2_X1 U728 ( .A(n814), .B(n1217), .Z(n1218) );
  INV_X4 U729 ( .A(in1[10]), .ZN(n976) );
  NOR2_X2 U730 ( .A1(n974), .A2(n977), .ZN(U8_Z_0) );
  INV_X4 U731 ( .A(in2[3]), .ZN(n978) );
  XNOR2_X2 U732 ( .A(U6_A_0_), .B(U6_B_0_), .ZN(n981) );
  NOR2_X2 U733 ( .A1(reset), .A2(n981), .ZN(U9_Z_0) );
  NOR2_X2 U734 ( .A1(n974), .A2(n984), .ZN(U8_Z_1) );
  NOR2_X2 U735 ( .A1(n974), .A2(n987), .ZN(U7_Z_1) );
  NAND2_X2 U736 ( .A1(U6_B_0_), .A2(U6_A_0_), .ZN(n1000) );
  NOR2_X2 U737 ( .A1(n974), .A2(n988), .ZN(U9_Z_1) );
  INV_X4 U738 ( .A(in3[1]), .ZN(n991) );
  OAI22_X2 U739 ( .A1(n778), .A2(n991), .B1(n989), .B2(n990), .ZN(n1005) );
  XNOR2_X2 U740 ( .A(net4221), .B(in1[12]), .ZN(n1007) );
  NOR2_X2 U741 ( .A1(n974), .A2(n992), .ZN(U8_Z_2) );
  INV_X4 U742 ( .A(in2[20]), .ZN(n1184) );
  NOR2_X2 U743 ( .A1(n973), .A2(n999), .ZN(U7_Z_2) );
  NOR2_X2 U744 ( .A1(U6_B_1_), .A2(U6_A_1_), .ZN(n1001) );
  NOR2_X2 U745 ( .A1(n973), .A2(n1004), .ZN(U9_Z_2) );
  INV_X4 U746 ( .A(in3[2]), .ZN(n1008) );
  OAI22_X2 U747 ( .A1(n1009), .A2(n1008), .B1(n1006), .B2(n1007), .ZN(n1023)
         );
  NOR2_X2 U748 ( .A1(n974), .A2(n1011), .ZN(U8_Z_3) );
  INV_X4 U749 ( .A(in2[21]), .ZN(n1196) );
  NOR2_X2 U750 ( .A1(n973), .A2(n1017), .ZN(U7_Z_3) );
  NOR2_X2 U751 ( .A1(U6_B_2_), .A2(U6_A_2_), .ZN(n1018) );
  OAI22_X2 U752 ( .A1(n1020), .A2(n1019), .B1(n927), .B2(n1018), .ZN(n1021) );
  NOR2_X2 U753 ( .A1(n974), .A2(n1022), .ZN(U9_Z_3) );
  INV_X4 U754 ( .A(in3[3]), .ZN(n1026) );
  OAI22_X2 U755 ( .A1(n1027), .A2(n1026), .B1(n1024), .B2(n1025), .ZN(n1038)
         );
  NOR2_X2 U756 ( .A1(n973), .A2(n1028), .ZN(U8_Z_4) );
  INV_X4 U757 ( .A(in2[22]), .ZN(n1206) );
  XOR2_X2 U758 ( .A(n1206), .B(in2[11]), .Z(n1033) );
  XOR2_X2 U759 ( .A(n1033), .B(n821), .Z(n1047) );
  NOR2_X2 U760 ( .A1(n974), .A2(n1035), .ZN(U7_Z_4) );
  NOR2_X2 U761 ( .A1(n973), .A2(n1037), .ZN(U9_Z_4) );
  INV_X4 U762 ( .A(in3[4]), .ZN(n1041) );
  OAI22_X2 U763 ( .A1(n1042), .A2(n1041), .B1(n1039), .B2(n1040), .ZN(n1056)
         );
  NOR2_X2 U764 ( .A1(n974), .A2(n1043), .ZN(U8_Z_5) );
  INV_X4 U765 ( .A(in2[23]), .ZN(n1224) );
  XOR2_X2 U766 ( .A(n1224), .B(in2[12]), .Z(n1048) );
  NOR2_X2 U767 ( .A1(reset), .A2(n1050), .ZN(U7_Z_5) );
  NOR2_X2 U768 ( .A1(U6_B_4_), .A2(U6_A_4_), .ZN(n1051) );
  OAI22_X2 U769 ( .A1(n1053), .A2(n1052), .B1(n924), .B2(n1051), .ZN(n1054) );
  NOR2_X2 U770 ( .A1(n973), .A2(n1055), .ZN(U9_Z_5) );
  NOR2_X2 U771 ( .A1(n1056), .A2(in3[5]), .ZN(n1057) );
  NOR2_X2 U772 ( .A1(n974), .A2(n1061), .ZN(U8_Z_6) );
  INV_X4 U773 ( .A(in2[24]), .ZN(n1237) );
  XOR2_X2 U774 ( .A(n1237), .B(in2[13]), .Z(n1065) );
  NOR2_X2 U775 ( .A1(n974), .A2(n1067), .ZN(U7_Z_6) );
  NOR2_X2 U776 ( .A1(n973), .A2(n1069), .ZN(U9_Z_6) );
  INV_X4 U777 ( .A(in3[6]), .ZN(n1073) );
  OAI22_X2 U778 ( .A1(n1074), .A2(n1073), .B1(n1071), .B2(n1072), .ZN(n1084)
         );
  XOR2_X2 U779 ( .A(in3[7]), .B(n932), .Z(n1075) );
  NOR2_X2 U780 ( .A1(n974), .A2(n1076), .ZN(U8_Z_7) );
  INV_X4 U781 ( .A(in2[25]), .ZN(n1251) );
  XOR2_X2 U782 ( .A(n1251), .B(in2[14]), .Z(n1077) );
  XOR2_X2 U783 ( .A(n1077), .B(in2[10]), .Z(n1091) );
  NOR2_X2 U784 ( .A1(n973), .A2(n1079), .ZN(U7_Z_7) );
  NOR2_X2 U785 ( .A1(U6_B_6_), .A2(U6_A_6_), .ZN(n1080) );
  NOR2_X2 U786 ( .A1(n974), .A2(n1083), .ZN(U9_Z_7) );
  NOR2_X2 U787 ( .A1(n974), .A2(n1087), .ZN(U8_Z_8) );
  NAND2_X2 U788 ( .A1(n1088), .A2(in4[7]), .ZN(n1089) );
  INV_X4 U789 ( .A(in2[26]), .ZN(n1263) );
  XOR2_X2 U790 ( .A(n1263), .B(in2[15]), .Z(n1092) );
  XOR2_X2 U791 ( .A(n1092), .B(in2[11]), .Z(n1105) );
  NOR2_X2 U792 ( .A1(n974), .A2(n1093), .ZN(U7_Z_8) );
  NOR2_X2 U793 ( .A1(U6_B_7_), .A2(U6_A_7_), .ZN(n1094) );
  NOR2_X2 U794 ( .A1(n974), .A2(n1097), .ZN(U9_Z_8) );
  INV_X4 U795 ( .A(in3[8]), .ZN(n1101) );
  OAI22_X2 U796 ( .A1(n772), .A2(n1101), .B1(n1099), .B2(n1100), .ZN(n1114) );
  XOR2_X2 U797 ( .A(net4044), .B(net4335), .Z(n1116) );
  NOR2_X2 U798 ( .A1(n974), .A2(n1102), .ZN(U8_Z_9) );
  INV_X4 U799 ( .A(in4[8]), .ZN(n1106) );
  OAI22_X2 U800 ( .A1(n1107), .A2(n1106), .B1(n1104), .B2(n1105), .ZN(n1121)
         );
  XOR2_X2 U801 ( .A(net4035), .B(in2[12]), .Z(n1122) );
  NOR2_X2 U802 ( .A1(n973), .A2(n1108), .ZN(U7_Z_9) );
  NOR2_X2 U803 ( .A1(U6_B_8_), .A2(U6_A_8_), .ZN(n1109) );
  OAI22_X2 U804 ( .A1(n1111), .A2(n1110), .B1(n921), .B2(n1109), .ZN(n1112) );
  NOR2_X2 U805 ( .A1(reset), .A2(n1113), .ZN(U9_Z_9) );
  INV_X4 U806 ( .A(in3[9]), .ZN(n1117) );
  OAI22_X2 U807 ( .A1(n1118), .A2(n1117), .B1(n1115), .B2(n1116), .ZN(net3999)
         );
  XOR2_X2 U808 ( .A(n1191), .B(in1[29]), .Z(n1119) );
  NOR2_X2 U809 ( .A1(n974), .A2(n1120), .ZN(U8_Z_10) );
  XOR2_X2 U810 ( .A(net4010), .B(in2[13]), .Z(n1128) );
  NOR2_X2 U811 ( .A1(reset), .A2(n1123), .ZN(U7_Z_10) );
  NOR2_X2 U812 ( .A1(n974), .A2(n1125), .ZN(U9_Z_10) );
  NOR2_X2 U813 ( .A1(n973), .A2(n1126), .ZN(U8_Z_11) );
  XOR2_X2 U814 ( .A(n1165), .B(in2[29]), .Z(n1130) );
  XOR2_X2 U815 ( .A(n1130), .B(in2[14]), .Z(n1140) );
  NOR2_X2 U816 ( .A1(n974), .A2(n1131), .ZN(U7_Z_11) );
  NOR2_X2 U817 ( .A1(U6_B_10_), .A2(U6_A_10_), .ZN(n1132) );
  OAI22_X2 U818 ( .A1(n1134), .A2(n1133), .B1(n915), .B2(n1132), .ZN(n1135) );
  NOR2_X2 U819 ( .A1(reset), .A2(n1136), .ZN(U9_Z_11) );
  INV_X4 U820 ( .A(in1[29]), .ZN(n1215) );
  XOR2_X2 U821 ( .A(n1215), .B(in1[31]), .Z(n1137) );
  XOR2_X2 U822 ( .A(n1137), .B(in1[22]), .Z(net3947) );
  NOR2_X2 U823 ( .A1(n973), .A2(n1138), .ZN(U8_Z_12) );
  INV_X4 U824 ( .A(in4[11]), .ZN(n1141) );
  OAI22_X2 U825 ( .A1(n835), .A2(n1141), .B1(n1139), .B2(n1140), .ZN(n1146) );
  XOR2_X2 U826 ( .A(n1148), .B(n1142), .Z(n1143) );
  NOR2_X2 U827 ( .A1(n974), .A2(n1143), .ZN(U7_Z_12) );
  NOR2_X2 U828 ( .A1(n973), .A2(n1145), .ZN(U9_Z_12) );
  NOR2_X2 U829 ( .A1(n974), .A2(net3941), .ZN(U8_Z_13) );
  NOR2_X2 U830 ( .A1(n974), .A2(n1150), .ZN(U7_Z_13) );
  NOR2_X2 U831 ( .A1(U6_B_12_), .A2(U6_A_12_), .ZN(n1151) );
  OAI22_X2 U832 ( .A1(n1153), .A2(n1152), .B1(n908), .B2(n1151), .ZN(n1154) );
  NOR2_X2 U833 ( .A1(n973), .A2(n1155), .ZN(U9_Z_13) );
  NOR2_X2 U834 ( .A1(n974), .A2(net3916), .ZN(U8_Z_14) );
  XOR2_X2 U835 ( .A(n1196), .B(in2[17]), .Z(n1164) );
  NOR2_X2 U836 ( .A1(n974), .A2(n1159), .ZN(U7_Z_14) );
  NOR2_X2 U837 ( .A1(n973), .A2(n1160), .ZN(U9_Z_14) );
  XOR2_X2 U838 ( .A(in3[15]), .B(in1[25]), .Z(n1161) );
  NOR2_X2 U839 ( .A1(n974), .A2(n1162), .ZN(U8_Z_15) );
  OAI22_X2 U840 ( .A1(n777), .A2(n656), .B1(n655), .B2(n1164), .ZN(n1174) );
  XOR2_X2 U841 ( .A(n1165), .B(in2[22]), .Z(n1176) );
  NOR2_X2 U842 ( .A1(n974), .A2(n1166), .ZN(U7_Z_15) );
  NOR2_X2 U843 ( .A1(U6_B_14_), .A2(U6_A_14_), .ZN(n1167) );
  OAI22_X2 U844 ( .A1(n1169), .A2(n1168), .B1(n909), .B2(n1167), .ZN(n1170) );
  NOR2_X2 U845 ( .A1(n974), .A2(n1171), .ZN(U9_Z_15) );
  NOR2_X2 U846 ( .A1(n973), .A2(n1173), .ZN(U8_Z_16) );
  XOR2_X2 U847 ( .A(n782), .B(in2[23]), .Z(n1182) );
  NOR2_X2 U848 ( .A1(n973), .A2(n1177), .ZN(U7_Z_16) );
  NOR2_X2 U849 ( .A1(n973), .A2(n1178), .ZN(U9_Z_16) );
  NOR2_X2 U850 ( .A1(n973), .A2(n1180), .ZN(U8_Z_17) );
  NOR2_X2 U851 ( .A1(n845), .A2(n830), .ZN(n1181) );
  XOR2_X2 U852 ( .A(n1184), .B(in2[24]), .Z(n1194) );
  NOR2_X2 U853 ( .A1(n973), .A2(n1185), .ZN(U7_Z_17) );
  NOR2_X2 U854 ( .A1(U6_B_16_), .A2(U6_A_16_), .ZN(n1186) );
  OAI22_X2 U855 ( .A1(n1188), .A2(n1187), .B1(n910), .B2(n1186), .ZN(n1189) );
  NOR2_X2 U856 ( .A1(n973), .A2(n1190), .ZN(U9_Z_17) );
  NOR2_X2 U857 ( .A1(n973), .A2(n1192), .ZN(U8_Z_18) );
  INV_X4 U858 ( .A(in4[17]), .ZN(n1195) );
  OAI22_X2 U859 ( .A1(n786), .A2(n1195), .B1(n1193), .B2(n1194), .ZN(n1201) );
  XOR2_X2 U860 ( .A(n1196), .B(in2[25]), .Z(n1203) );
  NOR2_X2 U861 ( .A1(n973), .A2(n1197), .ZN(U7_Z_18) );
  NOR2_X2 U862 ( .A1(n973), .A2(n1198), .ZN(U9_Z_18) );
  XOR2_X2 U863 ( .A(in3[19]), .B(in1[29]), .Z(n1199) );
  NOR2_X2 U864 ( .A1(n973), .A2(n1200), .ZN(U8_Z_19) );
  INV_X4 U865 ( .A(in4[18]), .ZN(n1204) );
  NOR2_X2 U866 ( .A1(n1201), .A2(in4[18]), .ZN(n1202) );
  OAI22_X2 U867 ( .A1(n1205), .A2(n1204), .B1(n1202), .B2(n1203), .ZN(n1219)
         );
  XOR2_X2 U868 ( .A(n1206), .B(in2[26]), .Z(n1221) );
  NOR2_X2 U869 ( .A1(n973), .A2(n1207), .ZN(U7_Z_19) );
  NOR2_X2 U870 ( .A1(U6_B_18_), .A2(U6_A_18_), .ZN(n1208) );
  OAI22_X2 U871 ( .A1(n1210), .A2(n1209), .B1(n916), .B2(n1208), .ZN(n1211) );
  NOR2_X2 U872 ( .A1(n973), .A2(n1212), .ZN(U9_Z_19) );
  INV_X4 U873 ( .A(in3[19]), .ZN(n1214) );
  NOR2_X2 U874 ( .A1(in3[19]), .A2(in1[29]), .ZN(n1213) );
  OAI22_X2 U875 ( .A1(n1215), .A2(n1214), .B1(n899), .B2(n1213), .ZN(n1216) );
  INV_X4 U876 ( .A(n1216), .ZN(n1228) );
  XOR2_X2 U877 ( .A(in3[20]), .B(in1[30]), .Z(n1217) );
  NOR2_X2 U878 ( .A1(n973), .A2(n1218), .ZN(U8_Z_20) );
  INV_X4 U879 ( .A(in4[19]), .ZN(n1222) );
  NOR2_X2 U880 ( .A1(n1219), .A2(in4[19]), .ZN(n1220) );
  OAI22_X2 U881 ( .A1(n1223), .A2(n1222), .B1(n1220), .B2(n1221), .ZN(n1232)
         );
  XOR2_X2 U882 ( .A(n1224), .B(in2[27]), .Z(n1234) );
  NOR2_X2 U883 ( .A1(n973), .A2(n1225), .ZN(U7_Z_20) );
  NOR2_X2 U884 ( .A1(n973), .A2(n1226), .ZN(U9_Z_20) );
  INV_X4 U885 ( .A(in3[20]), .ZN(n1229) );
  NOR2_X2 U886 ( .A1(in3[20]), .A2(in1[30]), .ZN(n1227) );
  NOR2_X2 U887 ( .A1(n974), .A2(n1231), .ZN(U8_Z_21) );
  INV_X4 U888 ( .A(in4[20]), .ZN(n1235) );
  NOR2_X2 U889 ( .A1(n1232), .A2(in4[20]), .ZN(n1233) );
  OAI22_X2 U890 ( .A1(n1236), .A2(n1235), .B1(n1233), .B2(n1234), .ZN(n1246)
         );
  XOR2_X2 U891 ( .A(n1237), .B(in2[28]), .Z(n1248) );
  NOR2_X2 U892 ( .A1(n973), .A2(n1238), .ZN(U7_Z_21) );
  NOR2_X2 U893 ( .A1(U6_B_20_), .A2(U6_A_20_), .ZN(n1239) );
  OAI22_X2 U894 ( .A1(n1241), .A2(n1240), .B1(n917), .B2(n1239), .ZN(n1242) );
  NOR2_X2 U895 ( .A1(reset), .A2(n1243), .ZN(U9_Z_21) );
  XOR2_X2 U896 ( .A(in3[22]), .B(in1[0]), .Z(n1244) );
  NOR2_X2 U897 ( .A1(n973), .A2(n1245), .ZN(U8_Z_22) );
  INV_X4 U898 ( .A(in4[21]), .ZN(n1249) );
  NOR2_X2 U899 ( .A1(n1246), .A2(in4[21]), .ZN(n1247) );
  OAI22_X2 U900 ( .A1(n1250), .A2(n1249), .B1(n1247), .B2(n1248), .ZN(n1259)
         );
  XOR2_X2 U901 ( .A(n1251), .B(in2[29]), .Z(n1261) );
  NOR2_X2 U902 ( .A1(n973), .A2(n1252), .ZN(U7_Z_22) );
  NOR2_X2 U903 ( .A1(n973), .A2(n1253), .ZN(U9_Z_22) );
  INV_X4 U904 ( .A(in1[0]), .ZN(n1256) );
  INV_X4 U905 ( .A(in3[22]), .ZN(n1255) );
  NOR2_X2 U906 ( .A1(in3[22]), .A2(in1[0]), .ZN(n1254) );
  OAI22_X2 U907 ( .A1(n1256), .A2(n1255), .B1(n900), .B2(n1254), .ZN(n1257) );
  NOR2_X2 U908 ( .A1(n974), .A2(n1258), .ZN(U8_Z_23) );
  XOR2_X2 U909 ( .A(n1263), .B(in2[30]), .Z(net3683) );
  NOR2_X2 U910 ( .A1(reset), .A2(n1264), .ZN(U7_Z_23) );
  NOR2_X2 U911 ( .A1(U6_B_22_), .A2(U6_A_22_), .ZN(n1265) );
  OAI22_X2 U912 ( .A1(n1267), .A2(n1266), .B1(n918), .B2(n1265), .ZN(n1268) );
  NOR2_X2 U913 ( .A1(n973), .A2(n1269), .ZN(U9_Z_23) );
  XOR2_X2 U914 ( .A(in3[24]), .B(in1[2]), .Z(n1271) );
  NOR2_X2 U915 ( .A1(reset), .A2(n1272), .ZN(U8_Z_24) );
  NOR2_X2 U916 ( .A1(n973), .A2(n1273), .ZN(U7_Z_24) );
  NOR2_X2 U917 ( .A1(n973), .A2(n1274), .ZN(U9_Z_24) );
  INV_X4 U918 ( .A(in1[2]), .ZN(n1277) );
  INV_X4 U919 ( .A(in3[24]), .ZN(n1276) );
  NOR2_X2 U920 ( .A1(in3[24]), .A2(in1[2]), .ZN(n1275) );
  OAI22_X2 U921 ( .A1(n1277), .A2(n1276), .B1(n904), .B2(n1275), .ZN(n1278) );
  INV_X4 U922 ( .A(n1278), .ZN(n1288) );
  NOR2_X2 U923 ( .A1(n973), .A2(n1279), .ZN(U8_Z_25) );
  NOR2_X2 U924 ( .A1(n973), .A2(n1281), .ZN(U7_Z_25) );
  NOR2_X2 U925 ( .A1(U6_B_24_), .A2(U6_A_24_), .ZN(n1282) );
  OAI22_X2 U926 ( .A1(n1284), .A2(n1283), .B1(n919), .B2(n1282), .ZN(n1285) );
  NOR2_X2 U927 ( .A1(n973), .A2(n1286), .ZN(U9_Z_25) );
  INV_X4 U928 ( .A(in1[3]), .ZN(n1290) );
  INV_X4 U929 ( .A(in3[25]), .ZN(n1289) );
  NOR2_X2 U930 ( .A1(in3[25]), .A2(in1[3]), .ZN(n1287) );
  OAI22_X2 U931 ( .A1(n1290), .A2(n1289), .B1(n1288), .B2(n1287), .ZN(n1291)
         );
  NOR2_X2 U932 ( .A1(n973), .A2(n1292), .ZN(U8_Z_26) );
  NAND2_X2 U933 ( .A1(in4[25]), .A2(in2[28]), .ZN(net3620) );
  NAND2_X2 U934 ( .A1(net3620), .A2(net3639), .ZN(n1293) );
  XNOR2_X2 U935 ( .A(net3637), .B(n1293), .ZN(n1294) );
  NOR2_X2 U936 ( .A1(n973), .A2(n1294), .ZN(U7_Z_26) );
  NOR2_X2 U937 ( .A1(n973), .A2(n1295), .ZN(U9_Z_26) );
  XOR2_X2 U938 ( .A(in3[27]), .B(in1[5]), .Z(n1296) );
  NOR2_X2 U939 ( .A1(n973), .A2(n1297), .ZN(U8_Z_27) );
  NOR2_X2 U940 ( .A1(n973), .A2(n1298), .ZN(U7_Z_27) );
  NOR2_X2 U941 ( .A1(U6_B_26_), .A2(U6_A_26_), .ZN(n1299) );
  OAI22_X2 U942 ( .A1(n1301), .A2(n1300), .B1(n920), .B2(n1299), .ZN(n1302) );
  NOR2_X2 U943 ( .A1(n973), .A2(n1303), .ZN(U9_Z_27) );
  XOR2_X2 U944 ( .A(in3[28]), .B(in1[6]), .Z(n1304) );
  NOR2_X2 U945 ( .A1(n973), .A2(n1305), .ZN(U8_Z_28) );
  NOR2_X2 U946 ( .A1(n974), .A2(n1306), .ZN(U7_Z_28) );
  NOR2_X2 U947 ( .A1(n974), .A2(n1307), .ZN(U9_Z_28) );
  XOR2_X2 U948 ( .A(in3[29]), .B(in1[7]), .Z(n1308) );
  INV_X4 U949 ( .A(in2[31]), .ZN(net3572) );
  INV_X4 U950 ( .A(in4[28]), .ZN(net3573) );
  NOR2_X2 U951 ( .A1(reset), .A2(n1310), .ZN(U7_Z_29) );
  NOR2_X2 U952 ( .A1(U6_B_28_), .A2(U6_A_28_), .ZN(n1311) );
  OAI22_X2 U953 ( .A1(n1313), .A2(n1312), .B1(n922), .B2(n1311), .ZN(n1314) );
  NOR2_X2 U954 ( .A1(reset), .A2(n1315), .ZN(U9_Z_29) );
  NOR2_X2 U955 ( .A1(n973), .A2(n1316), .ZN(U8_Z_30) );
  NAND2_X2 U956 ( .A1(net3548), .A2(n975), .ZN(n1317) );
  XOR2_X2 U957 ( .A(U6_B_30_), .B(U6_A_30_), .Z(n1318) );
  XOR2_X2 U958 ( .A(n926), .B(n1318), .Z(n1319) );
  NOR2_X2 U959 ( .A1(reset), .A2(n1319), .ZN(U9_Z_30) );
  NAND2_X2 U960 ( .A1(in4[30]), .A2(in2[1]), .ZN(net3525) );
  NAND2_X2 U961 ( .A1(net3523), .A2(n975), .ZN(net3512) );
  XNOR2_X2 U962 ( .A(U6_B_31_), .B(U6_A_31_), .ZN(n1324) );
  NOR2_X2 U963 ( .A1(U6_B_30_), .A2(U6_A_30_), .ZN(n1320) );
  OAI22_X2 U964 ( .A1(n1322), .A2(n1321), .B1(n926), .B2(n1320), .ZN(n1323) );
  XOR2_X2 U965 ( .A(n1324), .B(n1323), .Z(n1325) );
  NOR2_X2 U966 ( .A1(reset), .A2(n1325), .ZN(U9_Z_31) );
endmodule

