
module fp_2 ( clock, reset, in1, in2, in3, in4, ops_out );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  output [31:0] ops_out;
  input clock, reset;
  wire   U13_Z_0, U13_Z_1, U13_Z_2, U13_Z_3, U13_Z_4, U13_Z_5, U13_Z_6,
         U13_Z_7, U13_Z_8, U13_Z_9, U13_Z_10, U13_Z_11, U13_Z_12, U13_Z_13,
         U13_Z_14, U13_Z_15, U13_Z_16, U13_Z_17, U13_Z_18, U13_Z_19, U13_Z_20,
         U13_Z_21, U13_Z_22, U13_Z_23, U13_Z_24, U13_Z_25, U13_Z_26, U13_Z_27,
         U13_Z_28, U13_Z_29, U13_Z_30, U13_Z_31, U12_Z_0, U12_Z_1, U12_Z_2,
         U12_Z_3, U12_Z_4, U12_Z_5, U12_Z_6, U12_Z_7, U12_Z_8, U12_Z_9,
         U12_Z_10, U12_Z_11, U12_Z_12, U12_Z_13, U12_Z_14, U12_Z_15, U12_Z_16,
         U12_Z_17, U12_Z_18, U12_Z_19, U12_Z_20, U12_Z_21, U12_Z_22, U12_Z_23,
         U12_Z_24, U12_Z_25, U12_Z_26, U12_Z_27, U12_Z_28, U12_Z_29, U12_Z_30,
         U12_Z_31, U11_Z_0, U11_Z_1, U11_Z_2, U11_Z_3, U11_Z_4, U11_Z_5,
         U11_Z_6, U11_Z_7, U11_Z_8, U11_Z_9, U11_Z_10, U11_Z_11, U11_Z_12,
         U11_Z_13, U11_Z_14, U11_Z_22, U11_Z_23, U11_Z_24, U11_Z_25, U11_Z_26,
         U11_Z_27, U11_Z_28, U11_Z_29, U11_Z_30, U11_Z_31, U10_Z_0, U10_Z_1,
         U10_Z_2, U10_Z_3, U10_Z_4, U10_Z_5, U10_Z_6, U10_Z_7, U10_Z_8,
         U10_Z_9, U10_Z_10, U10_Z_11, U10_Z_12, U10_Z_13, U10_Z_14, U10_Z_15,
         U10_Z_16, U10_Z_17, U10_Z_18, U10_Z_19, U10_Z_20, U10_Z_21, U10_Z_22,
         U10_Z_23, U10_Z_24, U10_Z_29, U10_Z_30, U10_Z_31, U9_Z_0, U9_Z_1,
         U9_Z_2, U9_Z_3, U9_Z_4, U9_Z_5, U9_Z_6, U9_Z_7, U9_Z_8, U9_Z_9,
         U9_Z_10, U9_Z_11, U9_Z_12, U9_Z_13, U9_Z_14, U9_Z_15, U9_Z_16,
         U9_Z_17, U9_Z_18, U9_Z_19, U9_Z_20, U9_Z_21, U9_Z_22, U9_Z_23,
         U9_Z_24, U9_Z_25, U9_Z_26, U9_Z_27, U9_Z_28, U9_Z_29, U9_Z_30,
         U9_Z_31, U8_Z_0, U8_Z_1, U8_Z_2, U8_Z_3, U8_Z_4, U8_Z_5, U8_Z_6,
         U8_Z_7, U8_Z_8, U8_Z_9, U8_Z_10, U8_Z_11, U8_Z_12, U8_Z_13, U8_Z_14,
         U8_Z_15, U8_Z_16, U8_Z_17, U8_Z_18, U8_Z_19, U8_Z_20, U8_Z_21,
         U8_Z_22, U8_Z_23, U8_Z_24, U8_Z_25, U8_Z_26, U8_Z_27, U8_Z_28,
         U8_Z_29, U8_Z_30, U8_Z_31, U7_Z_0, U7_Z_1, U7_Z_2, U7_Z_3, U7_Z_4,
         U7_Z_5, U7_Z_6, U7_Z_7, U7_Z_8, U7_Z_9, U7_Z_10, U7_Z_11, U7_Z_12,
         U7_Z_13, U7_Z_14, U7_Z_15, U7_Z_16, U7_Z_17, U7_Z_18, U7_Z_19,
         U7_Z_20, U7_Z_21, U7_Z_22, U7_Z_23, U7_Z_24, U7_Z_25, U7_Z_26,
         U7_Z_27, U7_Z_28, U7_Z_29, U7_Z_30, U7_Z_31, U6_A_31_, U6_A_30_,
         U6_A_29_, U6_A_28_, U6_A_27_, U6_A_26_, U6_A_25_, U6_A_24_, U6_A_23_,
         U6_A_22_, U6_A_21_, U6_A_20_, U6_A_19_, U6_A_18_, U6_A_17_, U6_A_16_,
         U6_A_15_, U6_A_14_, U6_A_13_, U6_A_12_, U6_A_11_, U6_A_10_, U6_A_9_,
         U6_A_8_, U6_A_7_, U6_A_6_, U6_A_5_, U6_A_4_, U6_A_3_, U6_A_2_,
         U6_A_1_, U6_B_31_, U6_B_29_, U6_B_28_, U6_B_27_, U6_B_26_, U6_B_25_,
         U6_B_24_, U6_B_23_, U6_B_22_, U6_B_21_, U6_B_20_, U6_B_19_, U6_B_18_,
         U6_B_17_, U6_B_16_, U6_B_15_, U6_B_14_, U6_B_13_, U6_B_12_, U6_B_11_,
         U6_B_10_, U6_B_9_, U6_B_8_, U6_B_7_, U6_B_6_, U6_B_5_, U6_B_4_,
         U6_B_3_, U6_B_2_, U6_B_1_, U5_A_31_, U5_A_30_, U5_A_29_, U5_A_28_,
         U5_A_27_, U5_A_26_, U5_A_25_, U5_A_24_, U5_A_23_, U5_A_22_, U5_A_21_,
         U5_A_20_, U5_A_19_, U5_A_18_, U5_A_17_, U5_A_16_, U5_A_15_, U5_A_14_,
         U5_A_13_, U5_A_12_, U5_A_11_, U5_A_10_, U5_A_9_, U5_A_8_, U5_A_7_,
         U5_A_6_, U5_A_5_, U5_A_4_, U5_A_3_, U5_A_2_, U5_A_1_, U5_B_31_,
         U5_B_29_, U5_B_28_, U5_B_27_, U5_B_26_, U5_B_25_, U5_B_24_, U5_B_23_,
         U5_B_22_, U5_B_21_, U5_B_20_, U5_B_19_, U5_B_18_, U5_B_17_, U5_B_16_,
         U5_B_15_, U5_B_14_, U5_B_13_, U5_B_12_, U5_B_11_, U5_B_10_, U5_B_9_,
         U5_B_8_, U5_B_7_, U5_B_6_, U5_B_5_, U5_B_4_, U5_B_3_, U5_B_2_,
         U5_B_1_, U4_A_31_, U4_A_30_, U4_A_29_, U4_A_28_, U4_A_27_, U4_A_26_,
         U4_A_25_, U4_A_24_, U4_A_23_, U4_A_22_, U4_A_21_, U4_A_20_, U4_A_19_,
         U4_A_18_, U4_A_17_, U4_A_16_, U4_A_15_, U4_A_14_, U4_A_13_, U4_A_12_,
         U4_A_11_, U4_A_10_, U4_A_9_, U4_A_8_, U4_A_7_, U4_A_6_, U4_A_5_,
         U4_A_4_, U4_A_3_, U4_A_2_, U4_A_1_, U4_B_31_, U4_B_29_, U4_B_28_,
         U4_B_27_, U4_B_26_, U4_B_25_, U4_B_24_, U4_B_23_, U4_B_22_, U4_B_21_,
         U4_B_20_, U4_B_19_, U4_B_18_, U4_B_17_, U4_B_16_, U4_B_15_, U4_B_14_,
         U4_B_13_, U4_B_12_, U4_B_11_, U4_B_10_, U4_B_9_, U4_B_8_, U4_B_7_,
         U4_B_6_, U4_B_5_, U4_B_4_, U4_B_3_, U4_B_2_, U4_B_1_, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n771, n772, n773, n774,
         n775, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n812, n813, n814, n815, n816, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n853, n854, n855, n856, n857,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563;

  DFF_X1 in3_holding_reg_31_ ( .D(U13_Z_31), .CK(clock), .Q(U4_B_31_) );
  DFF_X2 in3_holding_reg_30_ ( .D(U13_Z_30), .CK(clock), .QN(n761) );
  DFF_X1 in3_holding_reg_29_ ( .D(U13_Z_29), .CK(clock), .Q(U4_B_29_) );
  DFF_X1 in3_holding_reg_28_ ( .D(U13_Z_28), .CK(clock), .Q(U4_B_28_), .QN(
        n1558) );
  DFF_X1 in3_holding_reg_27_ ( .D(U13_Z_27), .CK(clock), .Q(U4_B_27_), .QN(
        n765) );
  DFF_X1 in3_holding_reg_26_ ( .D(U13_Z_26), .CK(clock), .Q(U4_B_26_), .QN(
        n1557) );
  DFF_X1 in3_holding_reg_25_ ( .D(U13_Z_25), .CK(clock), .Q(U4_B_25_) );
  DFF_X1 in3_holding_reg_24_ ( .D(U13_Z_24), .CK(clock), .Q(U4_B_24_) );
  DFF_X1 in3_holding_reg_23_ ( .D(U13_Z_23), .CK(clock), .Q(U4_B_23_) );
  DFF_X1 in3_holding_reg_22_ ( .D(U13_Z_22), .CK(clock), .Q(U4_B_22_) );
  DFF_X1 in3_holding_reg_21_ ( .D(U13_Z_21), .CK(clock), .Q(U4_B_21_) );
  DFF_X1 in3_holding_reg_20_ ( .D(U13_Z_20), .CK(clock), .Q(U4_B_20_) );
  DFF_X1 in3_holding_reg_19_ ( .D(U13_Z_19), .CK(clock), .Q(U4_B_19_) );
  DFF_X1 in3_holding_reg_18_ ( .D(U13_Z_18), .CK(clock), .Q(U4_B_18_), .QN(
        n1539) );
  DFF_X1 in3_holding_reg_17_ ( .D(U13_Z_17), .CK(clock), .Q(U4_B_17_) );
  DFF_X1 in3_holding_reg_16_ ( .D(U13_Z_16), .CK(clock), .Q(U4_B_16_), .QN(
        n1517) );
  DFF_X1 in3_holding_reg_15_ ( .D(U13_Z_15), .CK(clock), .Q(U4_B_15_), .QN(
        n1505) );
  DFF_X1 in3_holding_reg_14_ ( .D(U13_Z_14), .CK(clock), .Q(U4_B_14_) );
  DFF_X1 in3_holding_reg_13_ ( .D(U13_Z_13), .CK(clock), .Q(U4_B_13_) );
  DFF_X1 in3_holding_reg_12_ ( .D(U13_Z_12), .CK(clock), .Q(U4_B_12_), .QN(
        n1537) );
  DFF_X1 in3_holding_reg_11_ ( .D(U13_Z_11), .CK(clock), .Q(U4_B_11_), .QN(
        n1534) );
  DFF_X1 in3_holding_reg_10_ ( .D(U13_Z_10), .CK(clock), .Q(U4_B_10_), .QN(
        n1514) );
  DFF_X1 in3_holding_reg_9_ ( .D(U13_Z_9), .CK(clock), .Q(U4_B_9_), .QN(n1499)
         );
  DFF_X1 in3_holding_reg_8_ ( .D(U13_Z_8), .CK(clock), .Q(U4_B_8_) );
  DFF_X1 in3_holding_reg_7_ ( .D(U13_Z_7), .CK(clock), .Q(U4_B_7_), .QN(n1555)
         );
  DFF_X1 in3_holding_reg_6_ ( .D(U13_Z_6), .CK(clock), .Q(U4_B_6_) );
  DFF_X1 in3_holding_reg_5_ ( .D(U13_Z_5), .CK(clock), .Q(U4_B_5_) );
  DFF_X1 in3_holding_reg_4_ ( .D(U13_Z_4), .CK(clock), .Q(U4_B_4_), .QN(n1533)
         );
  DFF_X1 in3_holding_reg_3_ ( .D(U13_Z_3), .CK(clock), .Q(U4_B_3_) );
  DFF_X1 in3_holding_reg_2_ ( .D(U13_Z_2), .CK(clock), .Q(U4_B_2_) );
  DFF_X1 in3_holding_reg_1_ ( .D(U13_Z_1), .CK(clock), .Q(U4_B_1_) );
  DFF_X2 in3_holding_reg_0_ ( .D(U13_Z_0), .CK(clock), .QN(n798) );
  DFF_X1 shift_1_reg_31_ ( .D(U11_Z_31), .CK(clock), .Q(U4_A_31_) );
  DFF_X1 shift_1_reg_30_ ( .D(U11_Z_30), .CK(clock), .Q(U4_A_30_), .QN(n799)
         );
  DFF_X1 shift_1_reg_29_ ( .D(U11_Z_29), .CK(clock), .Q(U4_A_29_) );
  DFF_X1 shift_1_reg_28_ ( .D(U11_Z_28), .CK(clock), .Q(U4_A_28_), .QN(n1559)
         );
  DFF_X1 shift_1_reg_27_ ( .D(U11_Z_27), .CK(clock), .Q(U4_A_27_), .QN(n800)
         );
  DFF_X1 shift_1_reg_26_ ( .D(U11_Z_26), .CK(clock), .Q(U4_A_26_), .QN(n1556)
         );
  DFF_X1 shift_1_reg_25_ ( .D(U11_Z_25), .CK(clock), .Q(U4_A_25_) );
  DFF_X1 shift_1_reg_24_ ( .D(U11_Z_24), .CK(clock), .Q(U4_A_24_) );
  DFF_X1 shift_1_reg_23_ ( .D(U11_Z_23), .CK(clock), .Q(U4_A_23_) );
  DFF_X1 shift_1_reg_22_ ( .D(U11_Z_22), .CK(clock), .Q(U4_A_22_) );
  SDFF_X1 shift_1_reg_21_ ( .D(in1[31]), .SI(1'b0), .SE(n1562), .CK(clock), 
        .Q(U4_A_21_) );
  SDFF_X1 shift_1_reg_20_ ( .D(in1[30]), .SI(1'b0), .SE(n1561), .CK(clock), 
        .Q(U4_A_20_) );
  SDFF_X1 shift_1_reg_19_ ( .D(in1[29]), .SI(1'b0), .SE(n1560), .CK(clock), 
        .Q(U4_A_19_) );
  SDFF_X1 shift_1_reg_18_ ( .D(in1[28]), .SI(1'b0), .SE(n1562), .CK(clock), 
        .Q(U4_A_18_), .QN(n1538) );
  SDFF_X1 shift_1_reg_17_ ( .D(in1[27]), .SI(1'b0), .SE(n1561), .CK(clock), 
        .Q(U4_A_17_) );
  SDFF_X1 shift_1_reg_16_ ( .D(in1[26]), .SI(1'b0), .SE(n1560), .CK(clock), 
        .Q(U4_A_16_), .QN(n1516) );
  SDFF_X1 shift_1_reg_15_ ( .D(in1[25]), .SI(1'b0), .SE(n1562), .CK(clock), 
        .Q(U4_A_15_), .QN(n1504) );
  DFF_X1 shift_1_reg_14_ ( .D(U11_Z_14), .CK(clock), .Q(U4_A_14_) );
  DFF_X1 shift_1_reg_13_ ( .D(U11_Z_13), .CK(clock), .Q(U4_A_13_) );
  DFF_X1 shift_1_reg_12_ ( .D(U11_Z_12), .CK(clock), .Q(U4_A_12_), .QN(n1536)
         );
  DFF_X1 shift_1_reg_11_ ( .D(U11_Z_11), .CK(clock), .Q(U4_A_11_), .QN(n1535)
         );
  DFF_X1 shift_1_reg_10_ ( .D(U11_Z_10), .CK(clock), .Q(U4_A_10_), .QN(n1515)
         );
  DFF_X1 shift_1_reg_9_ ( .D(U11_Z_9), .CK(clock), .Q(U4_A_9_), .QN(n1498) );
  DFF_X1 shift_1_reg_8_ ( .D(U11_Z_8), .CK(clock), .Q(U4_A_8_) );
  DFF_X1 shift_1_reg_7_ ( .D(U11_Z_7), .CK(clock), .Q(U4_A_7_), .QN(n1554) );
  DFF_X1 shift_1_reg_6_ ( .D(U11_Z_6), .CK(clock), .Q(U4_A_6_) );
  DFF_X1 shift_1_reg_5_ ( .D(U11_Z_5), .CK(clock), .Q(U4_A_5_) );
  DFF_X1 shift_1_reg_4_ ( .D(U11_Z_4), .CK(clock), .Q(U4_A_4_), .QN(n1532) );
  DFF_X1 shift_1_reg_3_ ( .D(U11_Z_3), .CK(clock), .Q(U4_A_3_) );
  DFF_X1 shift_1_reg_2_ ( .D(U11_Z_2), .CK(clock), .Q(U4_A_2_) );
  DFF_X1 shift_1_reg_1_ ( .D(U11_Z_1), .CK(clock), .Q(U4_A_1_) );
  DFF_X2 shift_1_reg_0_ ( .D(U11_Z_0), .CK(clock), .QN(n801) );
  DFF_X1 in4_holding_reg_31_ ( .D(U12_Z_31), .CK(clock), .Q(U5_B_31_) );
  DFF_X2 in4_holding_reg_30_ ( .D(U12_Z_30), .CK(clock), .QN(n802) );
  DFF_X1 in4_holding_reg_29_ ( .D(U12_Z_29), .CK(clock), .Q(U5_B_29_) );
  DFF_X1 in4_holding_reg_28_ ( .D(U12_Z_28), .CK(clock), .Q(U5_B_28_), .QN(
        n1552) );
  DFF_X1 in4_holding_reg_27_ ( .D(U12_Z_27), .CK(clock), .Q(U5_B_27_), .QN(
        n806) );
  DFF_X1 in4_holding_reg_26_ ( .D(U12_Z_26), .CK(clock), .Q(U5_B_26_), .QN(
        n1551) );
  DFF_X1 in4_holding_reg_25_ ( .D(U12_Z_25), .CK(clock), .Q(U5_B_25_) );
  DFF_X1 in4_holding_reg_24_ ( .D(U12_Z_24), .CK(clock), .Q(U5_B_24_) );
  DFF_X1 in4_holding_reg_23_ ( .D(U12_Z_23), .CK(clock), .Q(U5_B_23_) );
  DFF_X1 in4_holding_reg_22_ ( .D(U12_Z_22), .CK(clock), .Q(U5_B_22_) );
  DFF_X1 in4_holding_reg_21_ ( .D(U12_Z_21), .CK(clock), .Q(U5_B_21_) );
  DFF_X1 in4_holding_reg_20_ ( .D(U12_Z_20), .CK(clock), .Q(U5_B_20_) );
  DFF_X1 in4_holding_reg_19_ ( .D(U12_Z_19), .CK(clock), .Q(U5_B_19_) );
  DFF_X1 in4_holding_reg_18_ ( .D(U12_Z_18), .CK(clock), .Q(U5_B_18_), .QN(
        n1531) );
  DFF_X1 in4_holding_reg_17_ ( .D(U12_Z_17), .CK(clock), .Q(U5_B_17_) );
  DFF_X1 in4_holding_reg_16_ ( .D(U12_Z_16), .CK(clock), .Q(U5_B_16_), .QN(
        n1513) );
  DFF_X1 in4_holding_reg_15_ ( .D(U12_Z_15), .CK(clock), .Q(U5_B_15_), .QN(
        n1503) );
  DFF_X1 in4_holding_reg_14_ ( .D(U12_Z_14), .CK(clock), .Q(U5_B_14_) );
  DFF_X1 in4_holding_reg_13_ ( .D(U12_Z_13), .CK(clock), .Q(U5_B_13_) );
  DFF_X1 in4_holding_reg_12_ ( .D(U12_Z_12), .CK(clock), .Q(U5_B_12_), .QN(
        n1529) );
  DFF_X1 in4_holding_reg_11_ ( .D(U12_Z_11), .CK(clock), .Q(U5_B_11_), .QN(
        n1526) );
  DFF_X1 in4_holding_reg_10_ ( .D(U12_Z_10), .CK(clock), .Q(U5_B_10_), .QN(
        n1510) );
  DFF_X1 in4_holding_reg_9_ ( .D(U12_Z_9), .CK(clock), .Q(U5_B_9_), .QN(n1497)
         );
  DFF_X1 in4_holding_reg_8_ ( .D(U12_Z_8), .CK(clock), .Q(U5_B_8_) );
  DFF_X1 in4_holding_reg_7_ ( .D(U12_Z_7), .CK(clock), .Q(U5_B_7_), .QN(n1549)
         );
  DFF_X1 in4_holding_reg_6_ ( .D(U12_Z_6), .CK(clock), .Q(U5_B_6_) );
  DFF_X1 in4_holding_reg_5_ ( .D(U12_Z_5), .CK(clock), .Q(U5_B_5_) );
  DFF_X1 in4_holding_reg_4_ ( .D(U12_Z_4), .CK(clock), .Q(U5_B_4_), .QN(n1525)
         );
  DFF_X1 in4_holding_reg_3_ ( .D(U12_Z_3), .CK(clock), .Q(U5_B_3_) );
  DFF_X1 in4_holding_reg_2_ ( .D(U12_Z_2), .CK(clock), .Q(U5_B_2_) );
  DFF_X1 in4_holding_reg_1_ ( .D(U12_Z_1), .CK(clock), .Q(U5_B_1_) );
  DFF_X2 in4_holding_reg_0_ ( .D(U12_Z_0), .CK(clock), .QN(n839) );
  DFF_X1 shift_2_reg_31_ ( .D(U10_Z_31), .CK(clock), .Q(U5_A_31_) );
  DFF_X1 shift_2_reg_30_ ( .D(U10_Z_30), .CK(clock), .Q(U5_A_30_), .QN(n840)
         );
  DFF_X1 shift_2_reg_29_ ( .D(U10_Z_29), .CK(clock), .Q(U5_A_29_) );
  SDFF_X1 shift_2_reg_28_ ( .D(in2[31]), .SI(1'b0), .SE(n1561), .CK(clock), 
        .Q(U5_A_28_), .QN(n1553) );
  SDFF_X1 shift_2_reg_27_ ( .D(in2[30]), .SI(1'b0), .SE(n1560), .CK(clock), 
        .Q(U5_A_27_), .QN(n841) );
  SDFF_X1 shift_2_reg_26_ ( .D(in2[29]), .SI(1'b0), .SE(n1562), .CK(clock), 
        .Q(U5_A_26_), .QN(n1550) );
  SDFF_X1 shift_2_reg_25_ ( .D(in2[28]), .SI(1'b0), .SE(n1561), .CK(clock), 
        .Q(U5_A_25_) );
  DFF_X1 shift_2_reg_24_ ( .D(U10_Z_24), .CK(clock), .Q(U5_A_24_) );
  DFF_X1 shift_2_reg_23_ ( .D(U10_Z_23), .CK(clock), .Q(U5_A_23_) );
  DFF_X1 shift_2_reg_22_ ( .D(U10_Z_22), .CK(clock), .Q(U5_A_22_) );
  DFF_X1 shift_2_reg_21_ ( .D(U10_Z_21), .CK(clock), .Q(U5_A_21_) );
  DFF_X1 shift_2_reg_20_ ( .D(U10_Z_20), .CK(clock), .Q(U5_A_20_) );
  DFF_X1 shift_2_reg_19_ ( .D(U10_Z_19), .CK(clock), .Q(U5_A_19_) );
  DFF_X1 shift_2_reg_18_ ( .D(U10_Z_18), .CK(clock), .Q(U5_A_18_), .QN(n1530)
         );
  DFF_X1 shift_2_reg_17_ ( .D(U10_Z_17), .CK(clock), .Q(U5_A_17_) );
  DFF_X1 shift_2_reg_16_ ( .D(U10_Z_16), .CK(clock), .Q(U5_A_16_), .QN(n1512)
         );
  DFF_X1 shift_2_reg_15_ ( .D(U10_Z_15), .CK(clock), .Q(U5_A_15_), .QN(n1502)
         );
  DFF_X1 shift_2_reg_14_ ( .D(U10_Z_14), .CK(clock), .Q(U5_A_14_) );
  DFF_X1 shift_2_reg_13_ ( .D(U10_Z_13), .CK(clock), .Q(U5_A_13_) );
  DFF_X1 shift_2_reg_12_ ( .D(U10_Z_12), .CK(clock), .Q(U5_A_12_), .QN(n1528)
         );
  DFF_X1 shift_2_reg_11_ ( .D(U10_Z_11), .CK(clock), .Q(U5_A_11_), .QN(n1527)
         );
  DFF_X1 shift_2_reg_10_ ( .D(U10_Z_10), .CK(clock), .Q(U5_A_10_), .QN(n1511)
         );
  DFF_X1 shift_2_reg_9_ ( .D(U10_Z_9), .CK(clock), .Q(U5_A_9_), .QN(n1496) );
  DFF_X1 shift_2_reg_8_ ( .D(U10_Z_8), .CK(clock), .Q(U5_A_8_) );
  DFF_X1 shift_2_reg_7_ ( .D(U10_Z_7), .CK(clock), .Q(U5_A_7_), .QN(n1548) );
  DFF_X1 shift_2_reg_6_ ( .D(U10_Z_6), .CK(clock), .Q(U5_A_6_) );
  DFF_X1 shift_2_reg_5_ ( .D(U10_Z_5), .CK(clock), .Q(U5_A_5_) );
  DFF_X1 shift_2_reg_4_ ( .D(U10_Z_4), .CK(clock), .Q(U5_A_4_), .QN(n1524) );
  DFF_X1 shift_2_reg_3_ ( .D(U10_Z_3), .CK(clock), .Q(U5_A_3_) );
  DFF_X1 shift_2_reg_2_ ( .D(U10_Z_2), .CK(clock), .Q(U5_A_2_) );
  DFF_X1 shift_2_reg_1_ ( .D(U10_Z_1), .CK(clock), .Q(U5_A_1_) );
  DFF_X2 shift_2_reg_0_ ( .D(U10_Z_0), .CK(clock), .QN(n842) );
  DFF_X1 adr_1_op_reg_31_ ( .D(U8_Z_31), .CK(clock), .Q(U6_A_31_) );
  DFF_X1 adr_1_op_reg_30_ ( .D(U8_Z_30), .CK(clock), .Q(U6_A_30_), .QN(n843)
         );
  DFF_X1 adr_1_op_reg_29_ ( .D(U8_Z_29), .CK(clock), .Q(U6_A_29_) );
  DFF_X1 adr_1_op_reg_28_ ( .D(U8_Z_28), .CK(clock), .Q(U6_A_28_), .QN(n1521)
         );
  DFF_X1 adr_1_op_reg_27_ ( .D(U8_Z_27), .CK(clock), .Q(U6_A_27_), .QN(n847)
         );
  DFF_X1 adr_1_op_reg_26_ ( .D(U8_Z_26), .CK(clock), .Q(U6_A_26_), .QN(n1522)
         );
  DFF_X1 adr_1_op_reg_25_ ( .D(U8_Z_25), .CK(clock), .Q(U6_A_25_) );
  DFF_X1 adr_1_op_reg_24_ ( .D(U8_Z_24), .CK(clock), .Q(U6_A_24_) );
  DFF_X1 adr_1_op_reg_23_ ( .D(U8_Z_23), .CK(clock), .Q(U6_A_23_) );
  DFF_X1 adr_1_op_reg_22_ ( .D(U8_Z_22), .CK(clock), .Q(U6_A_22_) );
  DFF_X1 adr_1_op_reg_21_ ( .D(U8_Z_21), .CK(clock), .Q(U6_A_21_) );
  DFF_X1 adr_1_op_reg_20_ ( .D(U8_Z_20), .CK(clock), .Q(U6_A_20_) );
  DFF_X1 adr_1_op_reg_19_ ( .D(U8_Z_19), .CK(clock), .Q(U6_A_19_) );
  DFF_X1 adr_1_op_reg_18_ ( .D(U8_Z_18), .CK(clock), .Q(U6_A_18_), .QN(n1506)
         );
  DFF_X1 adr_1_op_reg_17_ ( .D(U8_Z_17), .CK(clock), .Q(U6_A_17_) );
  DFF_X1 adr_1_op_reg_16_ ( .D(U8_Z_16), .CK(clock), .Q(U6_A_16_), .QN(n1542)
         );
  DFF_X1 adr_1_op_reg_15_ ( .D(U8_Z_15), .CK(clock), .Q(U6_A_15_), .QN(n1500)
         );
  DFF_X1 adr_1_op_reg_14_ ( .D(U8_Z_14), .CK(clock), .Q(U6_A_14_) );
  DFF_X1 adr_1_op_reg_13_ ( .D(U8_Z_13), .CK(clock), .Q(U6_A_13_) );
  DFF_X1 adr_1_op_reg_12_ ( .D(U8_Z_12), .CK(clock), .Q(U6_A_12_), .QN(n1544)
         );
  DFF_X1 adr_1_op_reg_11_ ( .D(U8_Z_11), .CK(clock), .Q(U6_A_11_), .QN(n1495)
         );
  DFF_X1 adr_1_op_reg_10_ ( .D(U8_Z_10), .CK(clock), .Q(U6_A_10_), .QN(n1547)
         );
  DFF_X1 adr_1_op_reg_9_ ( .D(U8_Z_9), .CK(clock), .Q(U6_A_9_), .QN(n1508) );
  DFF_X1 adr_1_op_reg_8_ ( .D(U8_Z_8), .CK(clock), .Q(U6_A_8_) );
  DFF_X1 adr_1_op_reg_7_ ( .D(U8_Z_7), .CK(clock), .Q(U6_A_7_), .QN(n1518) );
  DFF_X1 adr_1_op_reg_6_ ( .D(U8_Z_6), .CK(clock), .Q(U6_A_6_) );
  DFF_X1 adr_1_op_reg_5_ ( .D(U8_Z_5), .CK(clock), .Q(U6_A_5_) );
  DFF_X1 adr_1_op_reg_4_ ( .D(U8_Z_4), .CK(clock), .Q(U6_A_4_), .QN(n1540) );
  DFF_X1 adr_1_op_reg_3_ ( .D(U8_Z_3), .CK(clock), .Q(U6_A_3_) );
  DFF_X1 adr_1_op_reg_2_ ( .D(U8_Z_2), .CK(clock), .Q(U6_A_2_) );
  DFF_X1 adr_1_op_reg_1_ ( .D(U8_Z_1), .CK(clock), .Q(U6_A_1_) );
  DFF_X2 adr_1_op_reg_0_ ( .D(U8_Z_0), .CK(clock), .QN(n880) );
  DFF_X1 adr_2_op_reg_31_ ( .D(U7_Z_31), .CK(clock), .Q(U6_B_31_) );
  DFF_X2 adr_2_op_reg_30_ ( .D(U7_Z_30), .CK(clock), .QN(n881) );
  DFF_X1 adr_2_op_reg_29_ ( .D(U7_Z_29), .CK(clock), .Q(U6_B_29_) );
  DFF_X1 adr_2_op_reg_28_ ( .D(U7_Z_28), .CK(clock), .Q(U6_B_28_), .QN(n1520)
         );
  DFF_X1 adr_2_op_reg_27_ ( .D(U7_Z_27), .CK(clock), .Q(U6_B_27_), .QN(n882)
         );
  DFF_X1 adr_2_op_reg_26_ ( .D(U7_Z_26), .CK(clock), .Q(U6_B_26_), .QN(n1523)
         );
  DFF_X1 adr_2_op_reg_25_ ( .D(U7_Z_25), .CK(clock), .Q(U6_B_25_) );
  DFF_X1 adr_2_op_reg_24_ ( .D(U7_Z_24), .CK(clock), .Q(U6_B_24_) );
  DFF_X1 adr_2_op_reg_23_ ( .D(U7_Z_23), .CK(clock), .Q(U6_B_23_) );
  DFF_X1 adr_2_op_reg_22_ ( .D(U7_Z_22), .CK(clock), .Q(U6_B_22_) );
  DFF_X1 adr_2_op_reg_21_ ( .D(U7_Z_21), .CK(clock), .Q(U6_B_21_) );
  DFF_X1 adr_2_op_reg_20_ ( .D(U7_Z_20), .CK(clock), .Q(U6_B_20_) );
  DFF_X1 adr_2_op_reg_19_ ( .D(U7_Z_19), .CK(clock), .Q(U6_B_19_) );
  DFF_X1 adr_2_op_reg_18_ ( .D(U7_Z_18), .CK(clock), .Q(U6_B_18_), .QN(n1507)
         );
  DFF_X1 adr_2_op_reg_17_ ( .D(U7_Z_17), .CK(clock), .Q(U6_B_17_) );
  DFF_X1 adr_2_op_reg_16_ ( .D(U7_Z_16), .CK(clock), .Q(U6_B_16_), .QN(n1543)
         );
  DFF_X1 adr_2_op_reg_15_ ( .D(U7_Z_15), .CK(clock), .Q(U6_B_15_), .QN(n1501)
         );
  DFF_X1 adr_2_op_reg_14_ ( .D(U7_Z_14), .CK(clock), .Q(U6_B_14_) );
  DFF_X1 adr_2_op_reg_13_ ( .D(U7_Z_13), .CK(clock), .Q(U6_B_13_) );
  DFF_X1 adr_2_op_reg_12_ ( .D(U7_Z_12), .CK(clock), .Q(U6_B_12_), .QN(n1545)
         );
  DFF_X1 adr_2_op_reg_11_ ( .D(U7_Z_11), .CK(clock), .Q(U6_B_11_), .QN(n1494)
         );
  DFF_X1 adr_2_op_reg_10_ ( .D(U7_Z_10), .CK(clock), .Q(U6_B_10_), .QN(n1546)
         );
  DFF_X1 adr_2_op_reg_9_ ( .D(U7_Z_9), .CK(clock), .Q(U6_B_9_), .QN(n1509) );
  DFF_X1 adr_2_op_reg_8_ ( .D(U7_Z_8), .CK(clock), .Q(U6_B_8_) );
  DFF_X1 adr_2_op_reg_7_ ( .D(U7_Z_7), .CK(clock), .Q(U6_B_7_), .QN(n1519) );
  DFF_X1 adr_2_op_reg_6_ ( .D(U7_Z_6), .CK(clock), .Q(U6_B_6_) );
  DFF_X1 adr_2_op_reg_5_ ( .D(U7_Z_5), .CK(clock), .Q(U6_B_5_) );
  DFF_X1 adr_2_op_reg_4_ ( .D(U7_Z_4), .CK(clock), .Q(U6_B_4_), .QN(n1541) );
  DFF_X1 adr_2_op_reg_3_ ( .D(U7_Z_3), .CK(clock), .Q(U6_B_3_) );
  DFF_X1 adr_2_op_reg_2_ ( .D(U7_Z_2), .CK(clock), .Q(U6_B_2_) );
  DFF_X1 adr_2_op_reg_1_ ( .D(U7_Z_1), .CK(clock), .Q(U6_B_1_) );
  DFF_X2 adr_2_op_reg_0_ ( .D(U7_Z_0), .CK(clock), .QN(n883) );
  NOR2_X2 U14 ( .A1(n1562), .A2(n890), .ZN(U9_Z_9) );
  XOR2_X2 U15 ( .A(n891), .B(n892), .Z(n890) );
  NOR2_X2 U18 ( .A1(n1560), .A2(n895), .ZN(U9_Z_8) );
  XOR2_X2 U19 ( .A(n893), .B(n896), .Z(n895) );
  NAND2_X2 U20 ( .A1(n872), .A2(n897), .ZN(n896) );
  NOR2_X2 U21 ( .A1(n1562), .A2(n899), .ZN(U9_Z_7) );
  XOR2_X2 U22 ( .A(n900), .B(n901), .Z(n899) );
  NOR2_X2 U24 ( .A1(n1561), .A2(n905), .ZN(U9_Z_6) );
  XOR2_X2 U25 ( .A(n904), .B(n906), .Z(n905) );
  NAND2_X2 U26 ( .A1(n874), .A2(n907), .ZN(n906) );
  NOR2_X2 U28 ( .A1(reset), .A2(n912), .ZN(U9_Z_5) );
  XNOR2_X2 U29 ( .A(n913), .B(n914), .ZN(n912) );
  NAND2_X2 U30 ( .A1(n915), .A2(n910), .ZN(n914) );
  NAND2_X2 U31 ( .A1(n916), .A2(n917), .ZN(n910) );
  NOR2_X2 U33 ( .A1(reset), .A2(n918), .ZN(U9_Z_4) );
  XOR2_X2 U34 ( .A(n916), .B(n919), .Z(n918) );
  NAND2_X2 U35 ( .A1(n915), .A2(n917), .ZN(n919) );
  NOR2_X2 U36 ( .A1(n1560), .A2(n920), .ZN(U9_Z_31) );
  XOR2_X2 U37 ( .A(n921), .B(n922), .Z(n920) );
  XNOR2_X2 U38 ( .A(U6_B_31_), .B(U6_A_31_), .ZN(n922) );
  OAI221_X2 U39 ( .B1(n923), .B2(n881), .C1(n924), .C2(n843), .A(n925), .ZN(
        n921) );
  NAND4_X2 U40 ( .A1(n926), .A2(n927), .A3(n845), .A4(n846), .ZN(n925) );
  NAND2_X2 U41 ( .A1(n843), .A2(n881), .ZN(n927) );
  NOR2_X2 U42 ( .A1(U6_A_30_), .A2(n844), .ZN(n923) );
  NOR2_X2 U43 ( .A1(n1561), .A2(n928), .ZN(U9_Z_30) );
  XOR2_X2 U44 ( .A(n929), .B(n930), .Z(n928) );
  XNOR2_X2 U45 ( .A(n881), .B(U6_A_30_), .ZN(n930) );
  NOR2_X2 U48 ( .A1(n934), .A2(n933), .ZN(n931) );
  NOR2_X2 U49 ( .A1(n1562), .A2(n935), .ZN(U9_Z_3) );
  XOR2_X2 U50 ( .A(n936), .B(n937), .Z(n935) );
  NAND2_X2 U51 ( .A1(n877), .A2(n938), .ZN(n937) );
  NOR2_X2 U53 ( .A1(U6_A_2_), .A2(U6_B_2_), .ZN(n940) );
  NOR2_X2 U54 ( .A1(n1561), .A2(n942), .ZN(U9_Z_29) );
  XOR2_X2 U55 ( .A(n943), .B(n944), .Z(n942) );
  NOR2_X2 U58 ( .A1(U6_B_29_), .A2(U6_A_29_), .ZN(n933) );
  NOR2_X2 U59 ( .A1(n1561), .A2(n945), .ZN(U9_Z_28) );
  XOR2_X2 U60 ( .A(n926), .B(n946), .Z(n945) );
  NOR2_X2 U61 ( .A1(U6_A_28_), .A2(U6_B_28_), .ZN(n934) );
  OAI221_X2 U62 ( .B1(n947), .B2(n882), .C1(n948), .C2(n847), .A(n949), .ZN(
        n926) );
  OAI221_X2 U63 ( .B1(U6_B_27_), .B2(U6_A_27_), .C1(n950), .C2(n849), .A(n951), 
        .ZN(n949) );
  NOR3_X2 U64 ( .A1(n953), .A2(n954), .A3(n955), .ZN(n950) );
  NOR2_X2 U65 ( .A1(n848), .A2(U6_A_27_), .ZN(n947) );
  NOR2_X2 U66 ( .A1(n1560), .A2(n956), .ZN(U9_Z_27) );
  XOR2_X2 U67 ( .A(n957), .B(n958), .Z(n956) );
  XNOR2_X2 U68 ( .A(n882), .B(U6_A_27_), .ZN(n958) );
  NOR2_X2 U70 ( .A1(n1560), .A2(n960), .ZN(U9_Z_26) );
  XOR2_X2 U71 ( .A(n959), .B(n961), .Z(n960) );
  NAND2_X2 U72 ( .A1(n951), .A2(n948), .ZN(n961) );
  NAND2_X2 U73 ( .A1(U6_B_26_), .A2(U6_A_26_), .ZN(n948) );
  NOR2_X2 U76 ( .A1(n1562), .A2(n963), .ZN(U9_Z_25) );
  XNOR2_X2 U77 ( .A(n964), .B(n965), .ZN(n963) );
  NOR2_X2 U80 ( .A1(U6_B_25_), .A2(U6_A_25_), .ZN(n955) );
  NOR2_X2 U81 ( .A1(n1562), .A2(n967), .ZN(U9_Z_24) );
  XOR2_X2 U82 ( .A(n953), .B(n968), .Z(n967) );
  NOR2_X2 U83 ( .A1(n954), .A2(n851), .ZN(n968) );
  NAND2_X2 U84 ( .A1(U6_B_24_), .A2(U6_A_24_), .ZN(n966) );
  NOR2_X2 U85 ( .A1(U6_A_24_), .A2(U6_B_24_), .ZN(n954) );
  AOI221_X2 U86 ( .B1(n969), .B2(U6_B_23_), .C1(n970), .C2(U6_A_23_), .A(n971), 
        .ZN(n953) );
  NOR4_X2 U87 ( .A1(n972), .A2(n973), .A3(n974), .A4(n975), .ZN(n971) );
  NOR2_X2 U90 ( .A1(n1561), .A2(n979), .ZN(U9_Z_23) );
  XNOR2_X2 U91 ( .A(n980), .B(n981), .ZN(n979) );
  XOR2_X2 U92 ( .A(U6_B_23_), .B(U6_A_23_), .Z(n981) );
  NOR2_X2 U94 ( .A1(n1561), .A2(n983), .ZN(U9_Z_22) );
  XNOR2_X2 U95 ( .A(n982), .B(n984), .ZN(n983) );
  NOR2_X2 U97 ( .A1(U6_A_22_), .A2(U6_B_22_), .ZN(n973) );
  NAND2_X2 U98 ( .A1(U6_B_22_), .A2(U6_A_22_), .ZN(n978) );
  NOR2_X2 U101 ( .A1(n1560), .A2(n986), .ZN(U9_Z_21) );
  XNOR2_X2 U102 ( .A(n987), .B(n988), .ZN(n986) );
  NOR2_X2 U105 ( .A1(U6_B_21_), .A2(U6_A_21_), .ZN(n974) );
  NOR2_X2 U106 ( .A1(n1560), .A2(n990), .ZN(U9_Z_20) );
  XOR2_X2 U107 ( .A(n976), .B(n991), .Z(n990) );
  NOR2_X2 U108 ( .A1(n972), .A2(n855), .ZN(n991) );
  NAND2_X2 U109 ( .A1(U6_B_20_), .A2(U6_A_20_), .ZN(n989) );
  NOR2_X2 U110 ( .A1(U6_A_20_), .A2(U6_B_20_), .ZN(n972) );
  OAI221_X2 U112 ( .B1(n995), .B2(n996), .C1(n997), .C2(n998), .A(n999), .ZN(
        n994) );
  NAND2_X2 U113 ( .A1(n1000), .A2(n857), .ZN(n998) );
  NOR2_X2 U114 ( .A1(n1562), .A2(n1002), .ZN(U9_Z_2) );
  XOR2_X2 U115 ( .A(n878), .B(n1003), .Z(n1002) );
  NOR2_X2 U117 ( .A1(n1562), .A2(n1004), .ZN(U9_Z_19) );
  XOR2_X2 U118 ( .A(n1005), .B(n1006), .Z(n1004) );
  NOR2_X2 U119 ( .A1(U6_A_19_), .A2(U6_B_19_), .ZN(n995) );
  NAND2_X2 U120 ( .A1(U6_B_19_), .A2(U6_A_19_), .ZN(n999) );
  AND3_X2 U122 ( .A1(n1000), .A2(n1007), .A3(n860), .ZN(n1001) );
  NOR2_X2 U123 ( .A1(n1561), .A2(n1008), .ZN(U9_Z_18) );
  XOR2_X2 U124 ( .A(n1009), .B(n1010), .Z(n1008) );
  NAND2_X2 U125 ( .A1(n996), .A2(n1000), .ZN(n1010) );
  NAND2_X2 U126 ( .A1(U6_B_18_), .A2(U6_A_18_), .ZN(n996) );
  NAND2_X2 U127 ( .A1(n997), .A2(n1011), .ZN(n1009) );
  NAND3_X2 U128 ( .A1(n1007), .A2(n992), .A3(n860), .ZN(n1011) );
  NOR2_X2 U130 ( .A1(n1561), .A2(n1013), .ZN(U9_Z_17) );
  XOR2_X2 U131 ( .A(n1014), .B(n1015), .Z(n1013) );
  NOR2_X2 U134 ( .A1(U6_B_17_), .A2(U6_A_17_), .ZN(n1012) );
  NOR2_X2 U135 ( .A1(n1560), .A2(n1017), .ZN(U9_Z_16) );
  XOR2_X2 U136 ( .A(n992), .B(n1018), .Z(n1017) );
  NAND2_X2 U137 ( .A1(n1007), .A2(n1016), .ZN(n1018) );
  NAND2_X2 U138 ( .A1(U6_B_16_), .A2(U6_A_16_), .ZN(n1016) );
  NAND4_X2 U142 ( .A1(n1028), .A2(n862), .A3(n893), .A4(n867), .ZN(n1021) );
  NAND4_X2 U143 ( .A1(n1029), .A2(n865), .A3(n1030), .A4(n863), .ZN(n1020) );
  NOR2_X2 U144 ( .A1(n1560), .A2(n1031), .ZN(U9_Z_15) );
  XOR2_X2 U145 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR2_X2 U146 ( .A(U6_B_15_), .B(U6_A_15_), .Z(n1033) );
  NOR2_X2 U148 ( .A1(n1562), .A2(n1035), .ZN(U9_Z_14) );
  XNOR2_X2 U149 ( .A(n1034), .B(n1036), .ZN(n1035) );
  NOR2_X2 U150 ( .A1(n864), .A2(n1025), .ZN(n1036) );
  NOR2_X2 U151 ( .A1(U6_A_14_), .A2(U6_B_14_), .ZN(n1025) );
  NAND2_X2 U152 ( .A1(U6_B_14_), .A2(U6_A_14_), .ZN(n1027) );
  NAND2_X2 U153 ( .A1(n1026), .A2(n1037), .ZN(n1034) );
  NAND3_X2 U154 ( .A1(n865), .A2(n1030), .A3(n1038), .ZN(n1037) );
  NOR2_X2 U156 ( .A1(n1561), .A2(n1040), .ZN(U9_Z_13) );
  XOR2_X2 U157 ( .A(n1041), .B(n1042), .Z(n1040) );
  NOR2_X2 U160 ( .A1(U6_B_13_), .A2(U6_A_13_), .ZN(n1039) );
  NOR2_X2 U161 ( .A1(n1562), .A2(n1044), .ZN(U9_Z_12) );
  XOR2_X2 U162 ( .A(n1038), .B(n1045), .Z(n1044) );
  NAND2_X2 U163 ( .A1(n1043), .A2(n1030), .ZN(n1045) );
  NAND2_X2 U164 ( .A1(U6_B_12_), .A2(U6_A_12_), .ZN(n1043) );
  NAND2_X2 U165 ( .A1(n1019), .A2(n1046), .ZN(n1038) );
  NAND3_X2 U166 ( .A1(n893), .A2(n867), .A3(n1028), .ZN(n1046) );
  AOI221_X2 U167 ( .B1(n867), .B2(n1047), .C1(n869), .C2(n1048), .A(n1049), 
        .ZN(n1019) );
  NOR2_X2 U168 ( .A1(n1050), .A2(n1051), .ZN(n1048) );
  NOR2_X2 U169 ( .A1(n1560), .A2(n1052), .ZN(U9_Z_11) );
  XOR2_X2 U170 ( .A(n1053), .B(n1054), .Z(n1052) );
  NOR2_X2 U171 ( .A1(n1049), .A2(n1051), .ZN(n1054) );
  NOR2_X2 U172 ( .A1(U6_A_11_), .A2(U6_B_11_), .ZN(n1051) );
  AOI221_X2 U173 ( .B1(n1028), .B2(n893), .C1(n869), .C2(n868), .A(n1047), 
        .ZN(n1053) );
  NOR3_X2 U174 ( .A1(n1050), .A2(n898), .A3(n894), .ZN(n1028) );
  NOR2_X2 U175 ( .A1(n1561), .A2(n1055), .ZN(U9_Z_10) );
  XOR2_X2 U176 ( .A(n1056), .B(n1057), .Z(n1055) );
  NOR2_X2 U177 ( .A1(n1050), .A2(n1047), .ZN(n1057) );
  NOR2_X2 U178 ( .A1(U6_A_10_), .A2(U6_B_10_), .ZN(n1050) );
  NAND2_X2 U181 ( .A1(U6_B_8_), .A2(U6_A_8_), .ZN(n897) );
  NAND2_X2 U182 ( .A1(n902), .A2(n1060), .ZN(n893) );
  NAND2_X2 U184 ( .A1(U6_B_6_), .A2(U6_A_6_), .ZN(n907) );
  NOR2_X2 U186 ( .A1(U6_B_6_), .A2(U6_A_6_), .ZN(n908) );
  NAND3_X2 U187 ( .A1(n917), .A2(n916), .A3(n875), .ZN(n1062) );
  NAND2_X2 U192 ( .A1(U6_B_3_), .A2(U6_A_3_), .ZN(n938) );
  NAND2_X2 U193 ( .A1(U6_B_2_), .A2(U6_A_2_), .ZN(n941) );
  NOR2_X2 U194 ( .A1(U6_A_3_), .A2(U6_B_3_), .ZN(n1063) );
  NAND2_X2 U196 ( .A1(U6_B_4_), .A2(U6_A_4_), .ZN(n915) );
  NOR2_X2 U197 ( .A1(U6_A_5_), .A2(U6_B_5_), .ZN(n909) );
  NAND2_X2 U198 ( .A1(U6_B_7_), .A2(U6_A_7_), .ZN(n902) );
  NOR2_X2 U199 ( .A1(n898), .A2(n894), .ZN(n1058) );
  NOR2_X2 U200 ( .A1(U6_B_9_), .A2(U6_A_9_), .ZN(n894) );
  NOR2_X2 U201 ( .A1(U6_A_8_), .A2(U6_B_8_), .ZN(n898) );
  NOR2_X2 U202 ( .A1(n1560), .A2(n1067), .ZN(U9_Z_1) );
  XNOR2_X2 U203 ( .A(n1065), .B(n1068), .ZN(n1067) );
  XOR2_X2 U204 ( .A(U6_B_1_), .B(U6_A_1_), .Z(n1068) );
  NOR2_X2 U206 ( .A1(n883), .A2(n880), .ZN(n1065) );
  NOR2_X2 U207 ( .A1(n1561), .A2(n1069), .ZN(U8_Z_9) );
  XOR2_X2 U208 ( .A(n1070), .B(n1071), .Z(n1069) );
  NOR2_X2 U211 ( .A1(n1560), .A2(n1074), .ZN(U8_Z_8) );
  XOR2_X2 U212 ( .A(n1072), .B(n1075), .Z(n1074) );
  NAND2_X2 U213 ( .A1(n790), .A2(n1076), .ZN(n1075) );
  NOR2_X2 U214 ( .A1(n1560), .A2(n1078), .ZN(U8_Z_7) );
  XOR2_X2 U215 ( .A(n1079), .B(n1080), .Z(n1078) );
  NOR2_X2 U217 ( .A1(n1562), .A2(n1084), .ZN(U8_Z_6) );
  XOR2_X2 U218 ( .A(n1083), .B(n1085), .Z(n1084) );
  NAND2_X2 U219 ( .A1(n792), .A2(n1086), .ZN(n1085) );
  NOR2_X2 U221 ( .A1(n1562), .A2(n1091), .ZN(U8_Z_5) );
  XNOR2_X2 U222 ( .A(n1092), .B(n1093), .ZN(n1091) );
  NAND2_X2 U223 ( .A1(n1094), .A2(n1089), .ZN(n1093) );
  NAND2_X2 U224 ( .A1(n1095), .A2(n1096), .ZN(n1089) );
  NOR2_X2 U226 ( .A1(n1561), .A2(n1097), .ZN(U8_Z_4) );
  XOR2_X2 U227 ( .A(n1095), .B(n1098), .Z(n1097) );
  NAND2_X2 U228 ( .A1(n1094), .A2(n1096), .ZN(n1098) );
  NOR2_X2 U229 ( .A1(n1561), .A2(n1099), .ZN(U8_Z_31) );
  XOR2_X2 U230 ( .A(n1100), .B(n1101), .Z(n1099) );
  XNOR2_X2 U231 ( .A(U4_B_31_), .B(U4_A_31_), .ZN(n1101) );
  OAI221_X2 U232 ( .B1(n1102), .B2(n761), .C1(n1103), .C2(n799), .A(n1104), 
        .ZN(n1100) );
  NAND4_X2 U233 ( .A1(n1105), .A2(n1106), .A3(n763), .A4(n764), .ZN(n1104) );
  NAND2_X2 U234 ( .A1(n799), .A2(n761), .ZN(n1106) );
  NOR2_X2 U235 ( .A1(U4_A_30_), .A2(n762), .ZN(n1102) );
  NOR2_X2 U236 ( .A1(n1560), .A2(n1107), .ZN(U8_Z_30) );
  XOR2_X2 U237 ( .A(n1108), .B(n1109), .Z(n1107) );
  XNOR2_X2 U238 ( .A(n761), .B(U4_A_30_), .ZN(n1109) );
  NOR2_X2 U241 ( .A1(n1113), .A2(n1112), .ZN(n1110) );
  NOR2_X2 U242 ( .A1(n1560), .A2(n1114), .ZN(U8_Z_3) );
  XOR2_X2 U243 ( .A(n1115), .B(n1116), .Z(n1114) );
  NAND2_X2 U244 ( .A1(n795), .A2(n1117), .ZN(n1116) );
  NOR2_X2 U246 ( .A1(U4_A_2_), .A2(U4_B_2_), .ZN(n1119) );
  NOR2_X2 U247 ( .A1(n1562), .A2(n1121), .ZN(U8_Z_29) );
  XOR2_X2 U248 ( .A(n1122), .B(n1123), .Z(n1121) );
  NOR2_X2 U251 ( .A1(U4_B_29_), .A2(U4_A_29_), .ZN(n1112) );
  NOR2_X2 U252 ( .A1(n1562), .A2(n1124), .ZN(U8_Z_28) );
  XOR2_X2 U253 ( .A(n1105), .B(n1125), .Z(n1124) );
  NOR2_X2 U254 ( .A1(U4_A_28_), .A2(U4_B_28_), .ZN(n1113) );
  OAI221_X2 U255 ( .B1(n1126), .B2(n765), .C1(n1127), .C2(n800), .A(n1128), 
        .ZN(n1105) );
  OAI221_X2 U256 ( .B1(U4_B_27_), .B2(U4_A_27_), .C1(n1129), .C2(n767), .A(
        n1130), .ZN(n1128) );
  NOR3_X2 U257 ( .A1(n1132), .A2(n1133), .A3(n1134), .ZN(n1129) );
  NOR2_X2 U258 ( .A1(n766), .A2(U4_A_27_), .ZN(n1126) );
  NOR2_X2 U259 ( .A1(n1561), .A2(n1135), .ZN(U8_Z_27) );
  XOR2_X2 U260 ( .A(n1136), .B(n1137), .Z(n1135) );
  XNOR2_X2 U261 ( .A(n765), .B(U4_A_27_), .ZN(n1137) );
  NOR2_X2 U263 ( .A1(n1561), .A2(n1139), .ZN(U8_Z_26) );
  XOR2_X2 U264 ( .A(n1138), .B(n1140), .Z(n1139) );
  NAND2_X2 U265 ( .A1(n1130), .A2(n1127), .ZN(n1140) );
  NAND2_X2 U266 ( .A1(U4_B_26_), .A2(U4_A_26_), .ZN(n1127) );
  NOR2_X2 U269 ( .A1(n1560), .A2(n1142), .ZN(U8_Z_25) );
  XNOR2_X2 U270 ( .A(n1143), .B(n1144), .ZN(n1142) );
  NOR2_X2 U273 ( .A1(U4_B_25_), .A2(U4_A_25_), .ZN(n1134) );
  NOR2_X2 U274 ( .A1(n1560), .A2(n1146), .ZN(U8_Z_24) );
  XOR2_X2 U275 ( .A(n1132), .B(n1147), .Z(n1146) );
  NOR2_X2 U276 ( .A1(n1133), .A2(n769), .ZN(n1147) );
  NAND2_X2 U277 ( .A1(U4_B_24_), .A2(U4_A_24_), .ZN(n1145) );
  NOR2_X2 U278 ( .A1(U4_A_24_), .A2(U4_B_24_), .ZN(n1133) );
  AOI221_X2 U279 ( .B1(n1148), .B2(U4_B_23_), .C1(n1149), .C2(U4_A_23_), .A(
        n1150), .ZN(n1132) );
  NOR4_X2 U280 ( .A1(n1151), .A2(n1152), .A3(n1153), .A4(n1154), .ZN(n1150) );
  NOR2_X2 U283 ( .A1(n1562), .A2(n1158), .ZN(U8_Z_23) );
  XNOR2_X2 U284 ( .A(n1159), .B(n1160), .ZN(n1158) );
  XOR2_X2 U285 ( .A(U4_B_23_), .B(U4_A_23_), .Z(n1160) );
  NOR2_X2 U287 ( .A1(n1562), .A2(n1162), .ZN(U8_Z_22) );
  XNOR2_X2 U288 ( .A(n1161), .B(n1163), .ZN(n1162) );
  NOR2_X2 U290 ( .A1(U4_A_22_), .A2(U4_B_22_), .ZN(n1152) );
  NAND2_X2 U291 ( .A1(U4_B_22_), .A2(U4_A_22_), .ZN(n1157) );
  NOR2_X2 U294 ( .A1(n1561), .A2(n1165), .ZN(U8_Z_21) );
  XNOR2_X2 U295 ( .A(n1166), .B(n1167), .ZN(n1165) );
  NOR2_X2 U298 ( .A1(U4_B_21_), .A2(U4_A_21_), .ZN(n1153) );
  NOR2_X2 U299 ( .A1(n1561), .A2(n1169), .ZN(U8_Z_20) );
  XOR2_X2 U300 ( .A(n1155), .B(n1170), .Z(n1169) );
  NOR2_X2 U301 ( .A1(n1151), .A2(n773), .ZN(n1170) );
  NAND2_X2 U302 ( .A1(U4_B_20_), .A2(U4_A_20_), .ZN(n1168) );
  NOR2_X2 U303 ( .A1(U4_A_20_), .A2(U4_B_20_), .ZN(n1151) );
  OAI221_X2 U305 ( .B1(n1174), .B2(n1175), .C1(n1176), .C2(n1177), .A(n1178), 
        .ZN(n1173) );
  NAND2_X2 U306 ( .A1(n1179), .A2(n775), .ZN(n1177) );
  NOR2_X2 U307 ( .A1(n1560), .A2(n1181), .ZN(U8_Z_2) );
  XOR2_X2 U308 ( .A(n796), .B(n1182), .Z(n1181) );
  NOR2_X2 U310 ( .A1(n1560), .A2(n1183), .ZN(U8_Z_19) );
  XOR2_X2 U311 ( .A(n1184), .B(n1185), .Z(n1183) );
  NOR2_X2 U312 ( .A1(U4_A_19_), .A2(U4_B_19_), .ZN(n1174) );
  NAND2_X2 U313 ( .A1(U4_B_19_), .A2(U4_A_19_), .ZN(n1178) );
  AND3_X2 U315 ( .A1(n1179), .A2(n1186), .A3(n778), .ZN(n1180) );
  NOR2_X2 U316 ( .A1(n1562), .A2(n1187), .ZN(U8_Z_18) );
  XOR2_X2 U317 ( .A(n1188), .B(n1189), .Z(n1187) );
  NAND2_X2 U318 ( .A1(n1175), .A2(n1179), .ZN(n1189) );
  NAND2_X2 U319 ( .A1(U4_B_18_), .A2(U4_A_18_), .ZN(n1175) );
  NAND2_X2 U320 ( .A1(n1176), .A2(n1190), .ZN(n1188) );
  NAND3_X2 U321 ( .A1(n1186), .A2(n1171), .A3(n778), .ZN(n1190) );
  NOR2_X2 U323 ( .A1(n1562), .A2(n1192), .ZN(U8_Z_17) );
  XOR2_X2 U324 ( .A(n1193), .B(n1194), .Z(n1192) );
  NOR2_X2 U327 ( .A1(U4_B_17_), .A2(U4_A_17_), .ZN(n1191) );
  NOR2_X2 U328 ( .A1(n1561), .A2(n1196), .ZN(U8_Z_16) );
  XOR2_X2 U329 ( .A(n1171), .B(n1197), .Z(n1196) );
  NAND2_X2 U330 ( .A1(n1186), .A2(n1195), .ZN(n1197) );
  NAND2_X2 U331 ( .A1(U4_B_16_), .A2(U4_A_16_), .ZN(n1195) );
  NAND4_X2 U335 ( .A1(n1207), .A2(n780), .A3(n1072), .A4(n785), .ZN(n1200) );
  NAND4_X2 U336 ( .A1(n1208), .A2(n783), .A3(n1209), .A4(n781), .ZN(n1199) );
  NOR2_X2 U337 ( .A1(n1561), .A2(n1210), .ZN(U8_Z_15) );
  XOR2_X2 U338 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR2_X2 U339 ( .A(U4_B_15_), .B(U4_A_15_), .Z(n1212) );
  NOR2_X2 U341 ( .A1(n1560), .A2(n1214), .ZN(U8_Z_14) );
  XNOR2_X2 U342 ( .A(n1213), .B(n1215), .ZN(n1214) );
  NOR2_X2 U343 ( .A1(n782), .A2(n1204), .ZN(n1215) );
  NOR2_X2 U344 ( .A1(U4_A_14_), .A2(U4_B_14_), .ZN(n1204) );
  NAND2_X2 U345 ( .A1(U4_B_14_), .A2(U4_A_14_), .ZN(n1206) );
  NAND2_X2 U346 ( .A1(n1205), .A2(n1216), .ZN(n1213) );
  NAND3_X2 U347 ( .A1(n783), .A2(n1209), .A3(n1217), .ZN(n1216) );
  NOR2_X2 U349 ( .A1(n1560), .A2(n1219), .ZN(U8_Z_13) );
  XOR2_X2 U350 ( .A(n1220), .B(n1221), .Z(n1219) );
  NOR2_X2 U353 ( .A1(U4_B_13_), .A2(U4_A_13_), .ZN(n1218) );
  NOR2_X2 U354 ( .A1(n1562), .A2(n1223), .ZN(U8_Z_12) );
  XOR2_X2 U355 ( .A(n1217), .B(n1224), .Z(n1223) );
  NAND2_X2 U356 ( .A1(n1222), .A2(n1209), .ZN(n1224) );
  NAND2_X2 U357 ( .A1(U4_B_12_), .A2(U4_A_12_), .ZN(n1222) );
  NAND2_X2 U358 ( .A1(n1198), .A2(n1225), .ZN(n1217) );
  NAND3_X2 U359 ( .A1(n1072), .A2(n785), .A3(n1207), .ZN(n1225) );
  AOI221_X2 U360 ( .B1(n785), .B2(n1226), .C1(n787), .C2(n1227), .A(n1228), 
        .ZN(n1198) );
  NOR2_X2 U361 ( .A1(n1229), .A2(n1230), .ZN(n1227) );
  NOR2_X2 U362 ( .A1(n1562), .A2(n1231), .ZN(U8_Z_11) );
  XOR2_X2 U363 ( .A(n1232), .B(n1233), .Z(n1231) );
  NOR2_X2 U364 ( .A1(n1228), .A2(n1230), .ZN(n1233) );
  NOR2_X2 U365 ( .A1(U4_A_11_), .A2(U4_B_11_), .ZN(n1230) );
  AOI221_X2 U366 ( .B1(n1207), .B2(n1072), .C1(n787), .C2(n786), .A(n1226), 
        .ZN(n1232) );
  NOR3_X2 U367 ( .A1(n1229), .A2(n1077), .A3(n1073), .ZN(n1207) );
  NOR2_X2 U368 ( .A1(n1561), .A2(n1234), .ZN(U8_Z_10) );
  XOR2_X2 U369 ( .A(n1235), .B(n1236), .Z(n1234) );
  NOR2_X2 U370 ( .A1(n1229), .A2(n1226), .ZN(n1236) );
  NOR2_X2 U371 ( .A1(U4_A_10_), .A2(U4_B_10_), .ZN(n1229) );
  NAND2_X2 U374 ( .A1(U4_B_8_), .A2(U4_A_8_), .ZN(n1076) );
  NAND2_X2 U375 ( .A1(n1081), .A2(n1239), .ZN(n1072) );
  NAND2_X2 U377 ( .A1(U4_B_6_), .A2(U4_A_6_), .ZN(n1086) );
  NOR2_X2 U379 ( .A1(U4_B_6_), .A2(U4_A_6_), .ZN(n1087) );
  NAND3_X2 U380 ( .A1(n1096), .A2(n1095), .A3(n793), .ZN(n1241) );
  NAND2_X2 U385 ( .A1(U4_B_3_), .A2(U4_A_3_), .ZN(n1117) );
  NAND2_X2 U386 ( .A1(U4_B_2_), .A2(U4_A_2_), .ZN(n1120) );
  NOR2_X2 U387 ( .A1(U4_A_3_), .A2(U4_B_3_), .ZN(n1242) );
  NAND2_X2 U389 ( .A1(U4_B_4_), .A2(U4_A_4_), .ZN(n1094) );
  NOR2_X2 U390 ( .A1(U4_A_5_), .A2(U4_B_5_), .ZN(n1088) );
  NAND2_X2 U391 ( .A1(U4_B_7_), .A2(U4_A_7_), .ZN(n1081) );
  NOR2_X2 U392 ( .A1(n1077), .A2(n1073), .ZN(n1237) );
  NOR2_X2 U393 ( .A1(U4_B_9_), .A2(U4_A_9_), .ZN(n1073) );
  NOR2_X2 U394 ( .A1(U4_A_8_), .A2(U4_B_8_), .ZN(n1077) );
  NOR2_X2 U395 ( .A1(n1561), .A2(n1246), .ZN(U8_Z_1) );
  XNOR2_X2 U396 ( .A(n1244), .B(n1247), .ZN(n1246) );
  XOR2_X2 U397 ( .A(U4_B_1_), .B(U4_A_1_), .Z(n1247) );
  NOR2_X2 U399 ( .A1(n798), .A2(n801), .ZN(n1244) );
  NOR2_X2 U400 ( .A1(n1560), .A2(n1248), .ZN(U7_Z_9) );
  XOR2_X2 U401 ( .A(n1249), .B(n1250), .Z(n1248) );
  NOR2_X2 U404 ( .A1(n1562), .A2(n1253), .ZN(U7_Z_8) );
  XOR2_X2 U405 ( .A(n1251), .B(n1254), .Z(n1253) );
  NAND2_X2 U406 ( .A1(n831), .A2(n1255), .ZN(n1254) );
  NOR2_X2 U407 ( .A1(n1561), .A2(n1257), .ZN(U7_Z_7) );
  XOR2_X2 U408 ( .A(n1258), .B(n1259), .Z(n1257) );
  NOR2_X2 U410 ( .A1(n1560), .A2(n1263), .ZN(U7_Z_6) );
  XOR2_X2 U411 ( .A(n1262), .B(n1264), .Z(n1263) );
  NAND2_X2 U412 ( .A1(n833), .A2(n1265), .ZN(n1264) );
  NOR2_X2 U414 ( .A1(n1562), .A2(n1270), .ZN(U7_Z_5) );
  XNOR2_X2 U415 ( .A(n1271), .B(n1272), .ZN(n1270) );
  NAND2_X2 U416 ( .A1(n1273), .A2(n1268), .ZN(n1272) );
  NAND2_X2 U417 ( .A1(n1274), .A2(n1275), .ZN(n1268) );
  NOR2_X2 U419 ( .A1(n1561), .A2(n1276), .ZN(U7_Z_4) );
  XOR2_X2 U420 ( .A(n1274), .B(n1277), .Z(n1276) );
  NAND2_X2 U421 ( .A1(n1273), .A2(n1275), .ZN(n1277) );
  NOR2_X2 U422 ( .A1(n1560), .A2(n1278), .ZN(U7_Z_31) );
  XOR2_X2 U423 ( .A(n1279), .B(n1280), .Z(n1278) );
  XNOR2_X2 U424 ( .A(U5_B_31_), .B(U5_A_31_), .ZN(n1280) );
  OAI221_X2 U425 ( .B1(n1281), .B2(n802), .C1(n1282), .C2(n840), .A(n1283), 
        .ZN(n1279) );
  NAND4_X2 U426 ( .A1(n1284), .A2(n1285), .A3(n804), .A4(n805), .ZN(n1283) );
  NAND2_X2 U427 ( .A1(n840), .A2(n802), .ZN(n1285) );
  NOR2_X2 U428 ( .A1(U5_A_30_), .A2(n803), .ZN(n1281) );
  NOR2_X2 U429 ( .A1(n1562), .A2(n1286), .ZN(U7_Z_30) );
  XOR2_X2 U430 ( .A(n1287), .B(n1288), .Z(n1286) );
  XNOR2_X2 U431 ( .A(n802), .B(U5_A_30_), .ZN(n1288) );
  NOR2_X2 U434 ( .A1(n1292), .A2(n1291), .ZN(n1289) );
  NOR2_X2 U435 ( .A1(n1562), .A2(n1293), .ZN(U7_Z_3) );
  XOR2_X2 U436 ( .A(n1294), .B(n1295), .Z(n1293) );
  NAND2_X2 U437 ( .A1(n836), .A2(n1296), .ZN(n1295) );
  NOR2_X2 U439 ( .A1(U5_A_2_), .A2(U5_B_2_), .ZN(n1298) );
  NOR2_X2 U440 ( .A1(n1561), .A2(n1300), .ZN(U7_Z_29) );
  XOR2_X2 U441 ( .A(n1301), .B(n1302), .Z(n1300) );
  NOR2_X2 U444 ( .A1(U5_B_29_), .A2(U5_A_29_), .ZN(n1291) );
  NOR2_X2 U445 ( .A1(n1560), .A2(n1303), .ZN(U7_Z_28) );
  XOR2_X2 U446 ( .A(n1284), .B(n1304), .Z(n1303) );
  NOR2_X2 U447 ( .A1(U5_A_28_), .A2(U5_B_28_), .ZN(n1292) );
  OAI221_X2 U448 ( .B1(n1305), .B2(n806), .C1(n1306), .C2(n841), .A(n1307), 
        .ZN(n1284) );
  OAI221_X2 U449 ( .B1(U5_B_27_), .B2(U5_A_27_), .C1(n1308), .C2(n808), .A(
        n1309), .ZN(n1307) );
  NOR3_X2 U450 ( .A1(n1311), .A2(n1312), .A3(n1313), .ZN(n1308) );
  NOR2_X2 U451 ( .A1(n807), .A2(U5_A_27_), .ZN(n1305) );
  NOR2_X2 U452 ( .A1(n1562), .A2(n1314), .ZN(U7_Z_27) );
  XOR2_X2 U453 ( .A(n1315), .B(n1316), .Z(n1314) );
  XNOR2_X2 U454 ( .A(n806), .B(U5_A_27_), .ZN(n1316) );
  NOR2_X2 U456 ( .A1(n1561), .A2(n1318), .ZN(U7_Z_26) );
  XOR2_X2 U457 ( .A(n1317), .B(n1319), .Z(n1318) );
  NAND2_X2 U458 ( .A1(n1309), .A2(n1306), .ZN(n1319) );
  NAND2_X2 U459 ( .A1(U5_B_26_), .A2(U5_A_26_), .ZN(n1306) );
  NOR2_X2 U462 ( .A1(n1560), .A2(n1321), .ZN(U7_Z_25) );
  XNOR2_X2 U463 ( .A(n1322), .B(n1323), .ZN(n1321) );
  NOR2_X2 U466 ( .A1(U5_B_25_), .A2(U5_A_25_), .ZN(n1313) );
  NOR2_X2 U467 ( .A1(n1562), .A2(n1325), .ZN(U7_Z_24) );
  XOR2_X2 U468 ( .A(n1311), .B(n1326), .Z(n1325) );
  NOR2_X2 U469 ( .A1(n1312), .A2(n810), .ZN(n1326) );
  NAND2_X2 U470 ( .A1(U5_B_24_), .A2(U5_A_24_), .ZN(n1324) );
  NOR2_X2 U471 ( .A1(U5_A_24_), .A2(U5_B_24_), .ZN(n1312) );
  AOI221_X2 U472 ( .B1(n1327), .B2(U5_B_23_), .C1(n1328), .C2(U5_A_23_), .A(
        n1329), .ZN(n1311) );
  NOR4_X2 U473 ( .A1(n1330), .A2(n1331), .A3(n1332), .A4(n1333), .ZN(n1329) );
  NOR2_X2 U476 ( .A1(n1561), .A2(n1337), .ZN(U7_Z_23) );
  XNOR2_X2 U477 ( .A(n1338), .B(n1339), .ZN(n1337) );
  XOR2_X2 U478 ( .A(U5_B_23_), .B(U5_A_23_), .Z(n1339) );
  NOR2_X2 U480 ( .A1(n1560), .A2(n1341), .ZN(U7_Z_22) );
  XNOR2_X2 U481 ( .A(n1340), .B(n1342), .ZN(n1341) );
  NOR2_X2 U483 ( .A1(U5_A_22_), .A2(U5_B_22_), .ZN(n1331) );
  NAND2_X2 U484 ( .A1(U5_B_22_), .A2(U5_A_22_), .ZN(n1336) );
  NOR2_X2 U487 ( .A1(n1562), .A2(n1344), .ZN(U7_Z_21) );
  XNOR2_X2 U488 ( .A(n1345), .B(n1346), .ZN(n1344) );
  NOR2_X2 U491 ( .A1(U5_B_21_), .A2(U5_A_21_), .ZN(n1332) );
  NOR2_X2 U492 ( .A1(n1561), .A2(n1348), .ZN(U7_Z_20) );
  XOR2_X2 U493 ( .A(n1334), .B(n1349), .Z(n1348) );
  NOR2_X2 U494 ( .A1(n1330), .A2(n814), .ZN(n1349) );
  NAND2_X2 U495 ( .A1(U5_B_20_), .A2(U5_A_20_), .ZN(n1347) );
  NOR2_X2 U496 ( .A1(U5_A_20_), .A2(U5_B_20_), .ZN(n1330) );
  OAI221_X2 U498 ( .B1(n1353), .B2(n1354), .C1(n1355), .C2(n1356), .A(n1357), 
        .ZN(n1352) );
  NAND2_X2 U499 ( .A1(n1358), .A2(n816), .ZN(n1356) );
  NOR2_X2 U500 ( .A1(n1560), .A2(n1360), .ZN(U7_Z_2) );
  XOR2_X2 U501 ( .A(n837), .B(n1361), .Z(n1360) );
  NOR2_X2 U503 ( .A1(n1562), .A2(n1362), .ZN(U7_Z_19) );
  XOR2_X2 U504 ( .A(n1363), .B(n1364), .Z(n1362) );
  NOR2_X2 U505 ( .A1(U5_A_19_), .A2(U5_B_19_), .ZN(n1353) );
  NAND2_X2 U506 ( .A1(U5_B_19_), .A2(U5_A_19_), .ZN(n1357) );
  AND3_X2 U508 ( .A1(n1358), .A2(n1365), .A3(n819), .ZN(n1359) );
  NOR2_X2 U509 ( .A1(n1561), .A2(n1366), .ZN(U7_Z_18) );
  XOR2_X2 U510 ( .A(n1367), .B(n1368), .Z(n1366) );
  NAND2_X2 U511 ( .A1(n1354), .A2(n1358), .ZN(n1368) );
  NAND2_X2 U512 ( .A1(U5_B_18_), .A2(U5_A_18_), .ZN(n1354) );
  NAND2_X2 U513 ( .A1(n1355), .A2(n1369), .ZN(n1367) );
  NAND3_X2 U514 ( .A1(n1365), .A2(n1350), .A3(n819), .ZN(n1369) );
  NOR2_X2 U516 ( .A1(n1560), .A2(n1371), .ZN(U7_Z_17) );
  XOR2_X2 U517 ( .A(n1372), .B(n1373), .Z(n1371) );
  NOR2_X2 U520 ( .A1(U5_B_17_), .A2(U5_A_17_), .ZN(n1370) );
  NOR2_X2 U521 ( .A1(n1562), .A2(n1375), .ZN(U7_Z_16) );
  XOR2_X2 U522 ( .A(n1350), .B(n1376), .Z(n1375) );
  NAND2_X2 U523 ( .A1(n1365), .A2(n1374), .ZN(n1376) );
  NAND2_X2 U524 ( .A1(U5_B_16_), .A2(U5_A_16_), .ZN(n1374) );
  NAND4_X2 U528 ( .A1(n1386), .A2(n821), .A3(n1251), .A4(n826), .ZN(n1379) );
  NAND4_X2 U529 ( .A1(n1387), .A2(n824), .A3(n1388), .A4(n822), .ZN(n1378) );
  NOR2_X2 U530 ( .A1(n1561), .A2(n1389), .ZN(U7_Z_15) );
  XOR2_X2 U531 ( .A(n1390), .B(n1391), .Z(n1389) );
  XOR2_X2 U532 ( .A(U5_B_15_), .B(U5_A_15_), .Z(n1391) );
  NOR2_X2 U534 ( .A1(n1560), .A2(n1393), .ZN(U7_Z_14) );
  XNOR2_X2 U535 ( .A(n1392), .B(n1394), .ZN(n1393) );
  NOR2_X2 U536 ( .A1(n823), .A2(n1383), .ZN(n1394) );
  NOR2_X2 U537 ( .A1(U5_A_14_), .A2(U5_B_14_), .ZN(n1383) );
  NAND2_X2 U538 ( .A1(U5_B_14_), .A2(U5_A_14_), .ZN(n1385) );
  NAND2_X2 U539 ( .A1(n1384), .A2(n1395), .ZN(n1392) );
  NAND3_X2 U540 ( .A1(n824), .A2(n1388), .A3(n1396), .ZN(n1395) );
  NOR2_X2 U542 ( .A1(n1562), .A2(n1398), .ZN(U7_Z_13) );
  XOR2_X2 U543 ( .A(n1399), .B(n1400), .Z(n1398) );
  NOR2_X2 U546 ( .A1(U5_B_13_), .A2(U5_A_13_), .ZN(n1397) );
  NOR2_X2 U547 ( .A1(n1560), .A2(n1402), .ZN(U7_Z_12) );
  XOR2_X2 U548 ( .A(n1396), .B(n1403), .Z(n1402) );
  NAND2_X2 U549 ( .A1(n1401), .A2(n1388), .ZN(n1403) );
  NAND2_X2 U550 ( .A1(U5_B_12_), .A2(U5_A_12_), .ZN(n1401) );
  NAND2_X2 U551 ( .A1(n1377), .A2(n1404), .ZN(n1396) );
  NAND3_X2 U552 ( .A1(n1251), .A2(n826), .A3(n1386), .ZN(n1404) );
  AOI221_X2 U553 ( .B1(n826), .B2(n1405), .C1(n828), .C2(n1406), .A(n1407), 
        .ZN(n1377) );
  NOR2_X2 U554 ( .A1(n1408), .A2(n1409), .ZN(n1406) );
  NOR2_X2 U555 ( .A1(n1562), .A2(n1410), .ZN(U7_Z_11) );
  XOR2_X2 U556 ( .A(n1411), .B(n1412), .Z(n1410) );
  NOR2_X2 U557 ( .A1(n1407), .A2(n1409), .ZN(n1412) );
  NOR2_X2 U558 ( .A1(U5_A_11_), .A2(U5_B_11_), .ZN(n1409) );
  AOI221_X2 U559 ( .B1(n1386), .B2(n1251), .C1(n828), .C2(n827), .A(n1405), 
        .ZN(n1411) );
  NOR3_X2 U560 ( .A1(n1408), .A2(n1256), .A3(n1252), .ZN(n1386) );
  NOR2_X2 U561 ( .A1(n1561), .A2(n1413), .ZN(U7_Z_10) );
  XOR2_X2 U562 ( .A(n1414), .B(n1415), .Z(n1413) );
  NOR2_X2 U563 ( .A1(n1408), .A2(n1405), .ZN(n1415) );
  NOR2_X2 U564 ( .A1(U5_A_10_), .A2(U5_B_10_), .ZN(n1408) );
  NAND2_X2 U567 ( .A1(U5_B_8_), .A2(U5_A_8_), .ZN(n1255) );
  NAND2_X2 U568 ( .A1(n1260), .A2(n1418), .ZN(n1251) );
  NAND2_X2 U570 ( .A1(U5_B_6_), .A2(U5_A_6_), .ZN(n1265) );
  NOR2_X2 U572 ( .A1(U5_B_6_), .A2(U5_A_6_), .ZN(n1266) );
  NAND3_X2 U573 ( .A1(n1275), .A2(n1274), .A3(n834), .ZN(n1420) );
  NAND2_X2 U578 ( .A1(U5_B_3_), .A2(U5_A_3_), .ZN(n1296) );
  NAND2_X2 U579 ( .A1(U5_B_2_), .A2(U5_A_2_), .ZN(n1299) );
  NOR2_X2 U580 ( .A1(U5_A_3_), .A2(U5_B_3_), .ZN(n1421) );
  NAND2_X2 U582 ( .A1(U5_B_4_), .A2(U5_A_4_), .ZN(n1273) );
  NOR2_X2 U583 ( .A1(U5_A_5_), .A2(U5_B_5_), .ZN(n1267) );
  NAND2_X2 U584 ( .A1(U5_B_7_), .A2(U5_A_7_), .ZN(n1260) );
  NOR2_X2 U585 ( .A1(n1256), .A2(n1252), .ZN(n1416) );
  NOR2_X2 U586 ( .A1(U5_B_9_), .A2(U5_A_9_), .ZN(n1252) );
  NOR2_X2 U587 ( .A1(U5_A_8_), .A2(U5_B_8_), .ZN(n1256) );
  NOR2_X2 U588 ( .A1(n1560), .A2(n1425), .ZN(U7_Z_1) );
  XNOR2_X2 U589 ( .A(n1423), .B(n1426), .ZN(n1425) );
  XOR2_X2 U590 ( .A(U5_B_1_), .B(U5_A_1_), .Z(n1426) );
  NOR2_X2 U592 ( .A1(n839), .A2(n842), .ZN(n1423) );
  NOR2_X2 U593 ( .A1(n1562), .A2(n1427), .ZN(U11_Z_9) );
  XNOR2_X2 U594 ( .A(in1[26]), .B(n1428), .ZN(n1427) );
  XOR2_X2 U595 ( .A(in1[19]), .B(in1[28]), .Z(n1428) );
  NOR2_X2 U596 ( .A1(n1561), .A2(n1429), .ZN(U11_Z_8) );
  XNOR2_X2 U597 ( .A(in1[25]), .B(n1430), .ZN(n1429) );
  XOR2_X2 U598 ( .A(in1[18]), .B(in1[27]), .Z(n1430) );
  NOR2_X2 U599 ( .A1(n1560), .A2(n1431), .ZN(U11_Z_7) );
  XNOR2_X2 U600 ( .A(in1[26]), .B(n1432), .ZN(n1431) );
  XOR2_X2 U601 ( .A(in1[24]), .B(in1[17]), .Z(n1432) );
  NOR2_X2 U602 ( .A1(n1562), .A2(n1433), .ZN(U11_Z_6) );
  XNOR2_X2 U603 ( .A(in1[25]), .B(n1434), .ZN(n1433) );
  XOR2_X2 U604 ( .A(in1[23]), .B(in1[16]), .Z(n1434) );
  NOR2_X2 U605 ( .A1(n1561), .A2(n1435), .ZN(U11_Z_5) );
  XOR2_X2 U606 ( .A(n1436), .B(in1[15]), .Z(n1435) );
  XNOR2_X2 U607 ( .A(in1[22]), .B(in1[24]), .ZN(n1436) );
  NOR2_X2 U608 ( .A1(n1560), .A2(n1437), .ZN(U11_Z_4) );
  XOR2_X2 U609 ( .A(n1438), .B(in1[14]), .Z(n1437) );
  XNOR2_X2 U610 ( .A(in1[21]), .B(in1[23]), .ZN(n1438) );
  NOR2_X2 U611 ( .A1(n1562), .A2(n1439), .ZN(U11_Z_3) );
  XOR2_X2 U612 ( .A(n1440), .B(in1[13]), .Z(n1439) );
  XNOR2_X2 U613 ( .A(in1[20]), .B(in1[22]), .ZN(n1440) );
  NOR2_X2 U614 ( .A1(n1561), .A2(n1441), .ZN(U11_Z_2) );
  XOR2_X2 U615 ( .A(n1442), .B(in1[12]), .Z(n1441) );
  XNOR2_X2 U616 ( .A(in1[19]), .B(in1[21]), .ZN(n1442) );
  NOR2_X2 U617 ( .A1(n1560), .A2(n1443), .ZN(U11_Z_14) );
  XNOR2_X2 U618 ( .A(in1[31]), .B(in1[24]), .ZN(n1443) );
  NOR2_X2 U619 ( .A1(n1562), .A2(n1444), .ZN(U11_Z_13) );
  XNOR2_X2 U620 ( .A(in1[30]), .B(in1[23]), .ZN(n1444) );
  NOR2_X2 U621 ( .A1(n1561), .A2(n1445), .ZN(U11_Z_12) );
  XNOR2_X2 U622 ( .A(in1[29]), .B(n1446), .ZN(n1445) );
  NOR2_X2 U624 ( .A1(n1560), .A2(n1447), .ZN(U11_Z_11) );
  XNOR2_X2 U625 ( .A(in1[28]), .B(n1448), .ZN(n1447) );
  NOR2_X2 U627 ( .A1(n1562), .A2(n1449), .ZN(U11_Z_10) );
  XNOR2_X2 U628 ( .A(in1[27]), .B(n1450), .ZN(n1449) );
  NOR2_X2 U630 ( .A1(n1561), .A2(n1451), .ZN(U11_Z_1) );
  XOR2_X2 U631 ( .A(n1452), .B(in1[11]), .Z(n1451) );
  XNOR2_X2 U632 ( .A(in1[18]), .B(in1[20]), .ZN(n1452) );
  NOR2_X2 U633 ( .A1(n1562), .A2(n1453), .ZN(U11_Z_0) );
  XOR2_X2 U634 ( .A(n1454), .B(in1[10]), .Z(n1453) );
  XNOR2_X2 U635 ( .A(in1[17]), .B(in1[19]), .ZN(n1454) );
  NOR2_X2 U636 ( .A1(n1560), .A2(n1455), .ZN(U10_Z_9) );
  XNOR2_X2 U637 ( .A(in2[12]), .B(n1456), .ZN(n1455) );
  XOR2_X2 U638 ( .A(in2[27]), .B(in2[16]), .Z(n1456) );
  NOR2_X2 U639 ( .A1(n1562), .A2(n1457), .ZN(U10_Z_8) );
  XNOR2_X2 U640 ( .A(in2[11]), .B(n1458), .ZN(n1457) );
  XOR2_X2 U641 ( .A(in2[26]), .B(in2[15]), .Z(n1458) );
  NOR2_X2 U642 ( .A1(n1561), .A2(n1459), .ZN(U10_Z_7) );
  XNOR2_X2 U643 ( .A(in2[10]), .B(n1460), .ZN(n1459) );
  XOR2_X2 U644 ( .A(in2[25]), .B(in2[14]), .Z(n1460) );
  NOR2_X2 U645 ( .A1(n1560), .A2(n1461), .ZN(U10_Z_6) );
  XNOR2_X2 U646 ( .A(in2[13]), .B(n1462), .ZN(n1461) );
  XOR2_X2 U647 ( .A(in2[9]), .B(in2[24]), .Z(n1462) );
  NOR2_X2 U648 ( .A1(n1562), .A2(n1463), .ZN(U10_Z_5) );
  XNOR2_X2 U649 ( .A(in2[12]), .B(n1464), .ZN(n1463) );
  XOR2_X2 U650 ( .A(in2[8]), .B(in2[23]), .Z(n1464) );
  NOR2_X2 U651 ( .A1(n1561), .A2(n1465), .ZN(U10_Z_4) );
  XNOR2_X2 U652 ( .A(in2[11]), .B(n1466), .ZN(n1465) );
  XOR2_X2 U653 ( .A(in2[7]), .B(in2[22]), .Z(n1466) );
  NOR2_X2 U654 ( .A1(n1560), .A2(n1467), .ZN(U10_Z_3) );
  XNOR2_X2 U655 ( .A(in2[10]), .B(n1468), .ZN(n1467) );
  XOR2_X2 U656 ( .A(in2[6]), .B(in2[21]), .Z(n1468) );
  NOR2_X2 U657 ( .A1(n1562), .A2(n1469), .ZN(U10_Z_24) );
  XNOR2_X2 U658 ( .A(in2[31]), .B(in2[27]), .ZN(n1469) );
  NOR2_X2 U659 ( .A1(n1561), .A2(n1470), .ZN(U10_Z_23) );
  XNOR2_X2 U660 ( .A(in2[30]), .B(in2[26]), .ZN(n1470) );
  NOR2_X2 U661 ( .A1(n1560), .A2(n1471), .ZN(U10_Z_22) );
  XNOR2_X2 U662 ( .A(in2[29]), .B(in2[25]), .ZN(n1471) );
  NOR2_X2 U663 ( .A1(n1561), .A2(n1472), .ZN(U10_Z_21) );
  XNOR2_X2 U664 ( .A(in2[28]), .B(in2[24]), .ZN(n1472) );
  NOR2_X2 U665 ( .A1(n1562), .A2(n1473), .ZN(U10_Z_20) );
  XNOR2_X2 U666 ( .A(in2[23]), .B(in2[27]), .ZN(n1473) );
  NOR2_X2 U667 ( .A1(n1560), .A2(n1474), .ZN(U10_Z_2) );
  XNOR2_X2 U668 ( .A(in2[20]), .B(n1475), .ZN(n1474) );
  XOR2_X2 U669 ( .A(in2[9]), .B(in2[5]), .Z(n1475) );
  NOR2_X2 U670 ( .A1(n1562), .A2(n1476), .ZN(U10_Z_19) );
  XNOR2_X2 U671 ( .A(in2[22]), .B(in2[26]), .ZN(n1476) );
  NOR2_X2 U672 ( .A1(n1561), .A2(n1477), .ZN(U10_Z_18) );
  XNOR2_X2 U673 ( .A(in2[21]), .B(in2[25]), .ZN(n1477) );
  NOR2_X2 U674 ( .A1(n1560), .A2(n1478), .ZN(U10_Z_17) );
  XNOR2_X2 U675 ( .A(in2[20]), .B(in2[24]), .ZN(n1478) );
  NOR2_X2 U676 ( .A1(n1562), .A2(n1479), .ZN(U10_Z_16) );
  XNOR2_X2 U677 ( .A(in2[19]), .B(in2[23]), .ZN(n1479) );
  NOR2_X2 U678 ( .A1(n1561), .A2(n1480), .ZN(U10_Z_15) );
  XNOR2_X2 U679 ( .A(in2[18]), .B(in2[22]), .ZN(n1480) );
  NOR2_X2 U680 ( .A1(n1560), .A2(n1481), .ZN(U10_Z_14) );
  XNOR2_X2 U681 ( .A(in2[17]), .B(in2[21]), .ZN(n1481) );
  NOR2_X2 U682 ( .A1(n1561), .A2(n1482), .ZN(U10_Z_13) );
  XNOR2_X2 U683 ( .A(in2[31]), .B(n1483), .ZN(n1482) );
  XOR2_X2 U684 ( .A(in2[20]), .B(in2[16]), .Z(n1483) );
  NOR2_X2 U685 ( .A1(n1560), .A2(n1484), .ZN(U10_Z_12) );
  XNOR2_X2 U686 ( .A(in2[30]), .B(n1485), .ZN(n1484) );
  NOR2_X2 U688 ( .A1(n1560), .A2(n1486), .ZN(U10_Z_11) );
  XNOR2_X2 U689 ( .A(in2[29]), .B(n1487), .ZN(n1486) );
  NOR2_X2 U691 ( .A1(n1562), .A2(n1488), .ZN(U10_Z_10) );
  XNOR2_X2 U692 ( .A(in2[28]), .B(n1489), .ZN(n1488) );
  XOR2_X2 U693 ( .A(in2[17]), .B(in2[13]), .Z(n1489) );
  NOR2_X2 U694 ( .A1(n1561), .A2(n1490), .ZN(U10_Z_1) );
  XNOR2_X2 U695 ( .A(in2[19]), .B(n1491), .ZN(n1490) );
  XOR2_X2 U696 ( .A(in2[8]), .B(in2[4]), .Z(n1491) );
  NOR2_X2 U697 ( .A1(n1560), .A2(n1492), .ZN(U10_Z_0) );
  XNOR2_X2 U698 ( .A(in2[18]), .B(n1493), .ZN(n1492) );
  XOR2_X2 U699 ( .A(in2[7]), .B(in2[3]), .Z(n1493) );
  INV_X4 U700 ( .A(n1103), .ZN(n762) );
  INV_X4 U701 ( .A(n1112), .ZN(n763) );
  INV_X4 U702 ( .A(n1113), .ZN(n764) );
  INV_X4 U703 ( .A(n1127), .ZN(n766) );
  INV_X4 U704 ( .A(n1131), .ZN(n767) );
  INV_X4 U705 ( .A(n1134), .ZN(n768) );
  INV_X4 U706 ( .A(n1145), .ZN(n769) );
  INV_X4 U708 ( .A(n1161), .ZN(n771) );
  INV_X4 U709 ( .A(n1153), .ZN(n772) );
  INV_X4 U710 ( .A(n1168), .ZN(n773) );
  INV_X4 U711 ( .A(n1155), .ZN(n774) );
  INV_X4 U712 ( .A(n1174), .ZN(n775) );
  INV_X4 U714 ( .A(n1176), .ZN(n777) );
  INV_X4 U715 ( .A(n1191), .ZN(n778) );
  INV_X4 U716 ( .A(n1195), .ZN(n779) );
  INV_X4 U717 ( .A(n1199), .ZN(n780) );
  INV_X4 U718 ( .A(n1204), .ZN(n781) );
  INV_X4 U719 ( .A(n1206), .ZN(n782) );
  INV_X4 U720 ( .A(n1218), .ZN(n783) );
  INV_X4 U721 ( .A(n1222), .ZN(n784) );
  INV_X4 U722 ( .A(n1230), .ZN(n785) );
  INV_X4 U723 ( .A(n1229), .ZN(n786) );
  INV_X4 U726 ( .A(n1076), .ZN(n789) );
  INV_X4 U727 ( .A(n1077), .ZN(n790) );
  INV_X4 U728 ( .A(n1086), .ZN(n791) );
  INV_X4 U729 ( .A(n1087), .ZN(n792) );
  INV_X4 U730 ( .A(n1088), .ZN(n793) );
  INV_X4 U731 ( .A(n1094), .ZN(n794) );
  INV_X4 U732 ( .A(n1242), .ZN(n795) );
  INV_X4 U733 ( .A(n1118), .ZN(n796) );
  INV_X4 U734 ( .A(n1245), .ZN(n797) );
  INV_X4 U735 ( .A(n1282), .ZN(n803) );
  INV_X4 U736 ( .A(n1291), .ZN(n804) );
  INV_X4 U737 ( .A(n1292), .ZN(n805) );
  INV_X4 U738 ( .A(n1306), .ZN(n807) );
  INV_X4 U739 ( .A(n1310), .ZN(n808) );
  INV_X4 U740 ( .A(n1313), .ZN(n809) );
  INV_X4 U741 ( .A(n1324), .ZN(n810) );
  INV_X4 U743 ( .A(n1340), .ZN(n812) );
  INV_X4 U744 ( .A(n1332), .ZN(n813) );
  INV_X4 U745 ( .A(n1347), .ZN(n814) );
  INV_X4 U746 ( .A(n1334), .ZN(n815) );
  INV_X4 U747 ( .A(n1353), .ZN(n816) );
  INV_X4 U749 ( .A(n1355), .ZN(n818) );
  INV_X4 U750 ( .A(n1370), .ZN(n819) );
  INV_X4 U751 ( .A(n1374), .ZN(n820) );
  INV_X4 U752 ( .A(n1378), .ZN(n821) );
  INV_X4 U753 ( .A(n1383), .ZN(n822) );
  INV_X4 U754 ( .A(n1385), .ZN(n823) );
  INV_X4 U755 ( .A(n1397), .ZN(n824) );
  INV_X4 U756 ( .A(n1401), .ZN(n825) );
  INV_X4 U757 ( .A(n1409), .ZN(n826) );
  INV_X4 U758 ( .A(n1408), .ZN(n827) );
  INV_X4 U761 ( .A(n1255), .ZN(n830) );
  INV_X4 U762 ( .A(n1256), .ZN(n831) );
  INV_X4 U763 ( .A(n1265), .ZN(n832) );
  INV_X4 U764 ( .A(n1266), .ZN(n833) );
  INV_X4 U765 ( .A(n1267), .ZN(n834) );
  INV_X4 U766 ( .A(n1273), .ZN(n835) );
  INV_X4 U767 ( .A(n1421), .ZN(n836) );
  INV_X4 U768 ( .A(n1297), .ZN(n837) );
  INV_X4 U769 ( .A(n1424), .ZN(n838) );
  INV_X4 U770 ( .A(n924), .ZN(n844) );
  INV_X4 U771 ( .A(n933), .ZN(n845) );
  INV_X4 U772 ( .A(n934), .ZN(n846) );
  INV_X4 U773 ( .A(n948), .ZN(n848) );
  INV_X4 U774 ( .A(n952), .ZN(n849) );
  INV_X4 U775 ( .A(n955), .ZN(n850) );
  INV_X4 U776 ( .A(n966), .ZN(n851) );
  INV_X4 U778 ( .A(n982), .ZN(n853) );
  INV_X4 U779 ( .A(n974), .ZN(n854) );
  INV_X4 U780 ( .A(n989), .ZN(n855) );
  INV_X4 U781 ( .A(n976), .ZN(n856) );
  INV_X4 U782 ( .A(n995), .ZN(n857) );
  INV_X4 U784 ( .A(n997), .ZN(n859) );
  INV_X4 U785 ( .A(n1012), .ZN(n860) );
  INV_X4 U786 ( .A(n1016), .ZN(n861) );
  INV_X4 U787 ( .A(n1020), .ZN(n862) );
  INV_X4 U788 ( .A(n1025), .ZN(n863) );
  INV_X4 U789 ( .A(n1027), .ZN(n864) );
  INV_X4 U790 ( .A(n1039), .ZN(n865) );
  INV_X4 U791 ( .A(n1043), .ZN(n866) );
  INV_X4 U792 ( .A(n1051), .ZN(n867) );
  INV_X4 U793 ( .A(n1050), .ZN(n868) );
  INV_X4 U796 ( .A(n897), .ZN(n871) );
  INV_X4 U797 ( .A(n898), .ZN(n872) );
  INV_X4 U798 ( .A(n907), .ZN(n873) );
  INV_X4 U799 ( .A(n908), .ZN(n874) );
  INV_X4 U800 ( .A(n909), .ZN(n875) );
  INV_X4 U801 ( .A(n915), .ZN(n876) );
  INV_X4 U802 ( .A(n1063), .ZN(n877) );
  INV_X4 U803 ( .A(n939), .ZN(n878) );
  INV_X4 U804 ( .A(n1066), .ZN(n879) );
  AND2_X1 U811 ( .A1(n902), .A2(n903), .ZN(n901) );
  OR2_X1 U812 ( .A1(n934), .A2(n932), .ZN(n946) );
  OR2_X1 U815 ( .A1(n955), .A2(n954), .ZN(n962) );
  OR2_X1 U816 ( .A1(U6_A_23_), .A2(n970), .ZN(n969) );
  OR2_X1 U817 ( .A1(n974), .A2(n972), .ZN(n985) );
  AND2_X1 U818 ( .A1(n1001), .A2(n857), .ZN(n993) );
  AND2_X1 U819 ( .A1(n999), .A2(n857), .ZN(n1006) );
  OR2_X1 U822 ( .A1(n1024), .A2(U6_A_15_), .ZN(n1023) );
  AND2_X1 U829 ( .A1(n1081), .A2(n1082), .ZN(n1080) );
  OR2_X1 U830 ( .A1(n1113), .A2(n1111), .ZN(n1125) );
  OR2_X1 U833 ( .A1(n1134), .A2(n1133), .ZN(n1141) );
  OR2_X1 U834 ( .A1(U4_A_23_), .A2(n1149), .ZN(n1148) );
  OR2_X1 U835 ( .A1(n1153), .A2(n1151), .ZN(n1164) );
  AND2_X1 U836 ( .A1(n1180), .A2(n775), .ZN(n1172) );
  AND2_X1 U837 ( .A1(n1178), .A2(n775), .ZN(n1185) );
  OR2_X1 U840 ( .A1(n1203), .A2(U4_A_15_), .ZN(n1202) );
  AND2_X1 U847 ( .A1(n1260), .A2(n1261), .ZN(n1259) );
  OR2_X1 U848 ( .A1(n1292), .A2(n1290), .ZN(n1304) );
  OR2_X1 U851 ( .A1(n1313), .A2(n1312), .ZN(n1320) );
  OR2_X1 U852 ( .A1(U5_A_23_), .A2(n1328), .ZN(n1327) );
  OR2_X1 U853 ( .A1(n1332), .A2(n1330), .ZN(n1343) );
  AND2_X1 U854 ( .A1(n1359), .A2(n816), .ZN(n1351) );
  AND2_X1 U855 ( .A1(n1357), .A2(n816), .ZN(n1364) );
  OR2_X1 U858 ( .A1(n1382), .A2(U5_A_15_), .ZN(n1381) );
  AND2_X1 U865 ( .A1(in3[9]), .A2(n1563), .ZN(U13_Z_9) );
  AND2_X1 U866 ( .A1(in3[8]), .A2(n1563), .ZN(U13_Z_8) );
  AND2_X1 U867 ( .A1(in3[7]), .A2(n1563), .ZN(U13_Z_7) );
  AND2_X1 U868 ( .A1(in3[6]), .A2(n1563), .ZN(U13_Z_6) );
  AND2_X1 U869 ( .A1(in3[5]), .A2(n1563), .ZN(U13_Z_5) );
  AND2_X1 U870 ( .A1(in3[4]), .A2(n1563), .ZN(U13_Z_4) );
  AND2_X1 U871 ( .A1(in3[31]), .A2(n1563), .ZN(U13_Z_31) );
  AND2_X1 U872 ( .A1(in3[30]), .A2(n1563), .ZN(U13_Z_30) );
  AND2_X1 U873 ( .A1(in3[3]), .A2(n1563), .ZN(U13_Z_3) );
  AND2_X1 U874 ( .A1(in3[29]), .A2(n1563), .ZN(U13_Z_29) );
  AND2_X1 U875 ( .A1(in3[28]), .A2(n1563), .ZN(U13_Z_28) );
  AND2_X1 U876 ( .A1(in3[27]), .A2(n1563), .ZN(U13_Z_27) );
  AND2_X1 U877 ( .A1(in3[26]), .A2(n1563), .ZN(U13_Z_26) );
  AND2_X1 U878 ( .A1(in3[25]), .A2(n1563), .ZN(U13_Z_25) );
  AND2_X1 U879 ( .A1(in3[24]), .A2(n1563), .ZN(U13_Z_24) );
  AND2_X1 U880 ( .A1(in3[23]), .A2(n1563), .ZN(U13_Z_23) );
  AND2_X1 U881 ( .A1(in3[22]), .A2(n1563), .ZN(U13_Z_22) );
  AND2_X1 U882 ( .A1(in3[21]), .A2(n1563), .ZN(U13_Z_21) );
  AND2_X1 U883 ( .A1(in3[20]), .A2(n1563), .ZN(U13_Z_20) );
  AND2_X1 U884 ( .A1(in3[2]), .A2(n1563), .ZN(U13_Z_2) );
  AND2_X1 U885 ( .A1(in3[19]), .A2(n1563), .ZN(U13_Z_19) );
  AND2_X1 U886 ( .A1(in3[18]), .A2(n1563), .ZN(U13_Z_18) );
  AND2_X1 U887 ( .A1(in3[17]), .A2(n1563), .ZN(U13_Z_17) );
  AND2_X1 U888 ( .A1(in3[16]), .A2(n1563), .ZN(U13_Z_16) );
  AND2_X1 U889 ( .A1(in3[15]), .A2(n1563), .ZN(U13_Z_15) );
  AND2_X1 U890 ( .A1(in3[14]), .A2(n1563), .ZN(U13_Z_14) );
  AND2_X1 U891 ( .A1(in3[13]), .A2(n1563), .ZN(U13_Z_13) );
  AND2_X1 U892 ( .A1(in3[12]), .A2(n1563), .ZN(U13_Z_12) );
  AND2_X1 U893 ( .A1(in3[11]), .A2(n1563), .ZN(U13_Z_11) );
  AND2_X1 U894 ( .A1(in3[10]), .A2(n1563), .ZN(U13_Z_10) );
  AND2_X1 U895 ( .A1(in3[1]), .A2(n1563), .ZN(U13_Z_1) );
  AND2_X1 U896 ( .A1(in3[0]), .A2(n1563), .ZN(U13_Z_0) );
  AND2_X1 U897 ( .A1(in4[9]), .A2(n1563), .ZN(U12_Z_9) );
  AND2_X1 U898 ( .A1(in4[8]), .A2(n1563), .ZN(U12_Z_8) );
  AND2_X1 U899 ( .A1(in4[7]), .A2(n1563), .ZN(U12_Z_7) );
  AND2_X1 U900 ( .A1(in4[6]), .A2(n1563), .ZN(U12_Z_6) );
  AND2_X1 U901 ( .A1(in4[5]), .A2(n1563), .ZN(U12_Z_5) );
  AND2_X1 U902 ( .A1(in4[4]), .A2(n1563), .ZN(U12_Z_4) );
  AND2_X1 U903 ( .A1(in4[31]), .A2(n1563), .ZN(U12_Z_31) );
  AND2_X1 U904 ( .A1(in4[30]), .A2(n1563), .ZN(U12_Z_30) );
  AND2_X1 U905 ( .A1(in4[3]), .A2(n1563), .ZN(U12_Z_3) );
  AND2_X1 U906 ( .A1(in4[29]), .A2(n1563), .ZN(U12_Z_29) );
  AND2_X1 U907 ( .A1(in4[28]), .A2(n1563), .ZN(U12_Z_28) );
  AND2_X1 U908 ( .A1(in4[27]), .A2(n1563), .ZN(U12_Z_27) );
  AND2_X1 U909 ( .A1(in4[26]), .A2(n1563), .ZN(U12_Z_26) );
  AND2_X1 U910 ( .A1(in4[25]), .A2(n1563), .ZN(U12_Z_25) );
  AND2_X1 U911 ( .A1(in4[24]), .A2(n1563), .ZN(U12_Z_24) );
  AND2_X1 U912 ( .A1(in4[23]), .A2(n1563), .ZN(U12_Z_23) );
  AND2_X1 U913 ( .A1(in4[22]), .A2(n1563), .ZN(U12_Z_22) );
  AND2_X1 U914 ( .A1(in4[21]), .A2(n1563), .ZN(U12_Z_21) );
  AND2_X1 U915 ( .A1(in4[20]), .A2(n1563), .ZN(U12_Z_20) );
  AND2_X1 U916 ( .A1(in4[2]), .A2(n1563), .ZN(U12_Z_2) );
  AND2_X1 U917 ( .A1(in4[19]), .A2(n1563), .ZN(U12_Z_19) );
  AND2_X1 U918 ( .A1(in4[18]), .A2(n1563), .ZN(U12_Z_18) );
  AND2_X1 U919 ( .A1(in4[17]), .A2(n1563), .ZN(U12_Z_17) );
  AND2_X1 U920 ( .A1(in4[16]), .A2(n1563), .ZN(U12_Z_16) );
  AND2_X1 U921 ( .A1(in4[15]), .A2(n1563), .ZN(U12_Z_15) );
  AND2_X1 U922 ( .A1(in4[14]), .A2(n1563), .ZN(U12_Z_14) );
  AND2_X1 U923 ( .A1(in4[13]), .A2(n1563), .ZN(U12_Z_13) );
  AND2_X1 U924 ( .A1(in4[12]), .A2(n1563), .ZN(U12_Z_12) );
  AND2_X1 U925 ( .A1(in4[11]), .A2(n1563), .ZN(U12_Z_11) );
  AND2_X1 U926 ( .A1(in4[10]), .A2(n1563), .ZN(U12_Z_10) );
  AND2_X1 U927 ( .A1(in4[1]), .A2(n1563), .ZN(U12_Z_1) );
  AND2_X1 U928 ( .A1(in4[0]), .A2(n1563), .ZN(U12_Z_0) );
  AND2_X1 U929 ( .A1(in1[9]), .A2(n1563), .ZN(U11_Z_31) );
  AND2_X1 U930 ( .A1(in1[8]), .A2(n1563), .ZN(U11_Z_30) );
  AND2_X1 U931 ( .A1(in1[7]), .A2(n1563), .ZN(U11_Z_29) );
  AND2_X1 U932 ( .A1(in1[6]), .A2(n1563), .ZN(U11_Z_28) );
  AND2_X1 U933 ( .A1(in1[5]), .A2(n1563), .ZN(U11_Z_27) );
  AND2_X1 U934 ( .A1(in1[4]), .A2(n1563), .ZN(U11_Z_26) );
  AND2_X1 U935 ( .A1(in1[3]), .A2(n1563), .ZN(U11_Z_25) );
  AND2_X1 U936 ( .A1(in1[2]), .A2(n1563), .ZN(U11_Z_24) );
  AND2_X1 U937 ( .A1(in1[1]), .A2(n1563), .ZN(U11_Z_23) );
  AND2_X1 U938 ( .A1(in1[0]), .A2(n1563), .ZN(U11_Z_22) );
  AND2_X1 U939 ( .A1(in2[2]), .A2(n1563), .ZN(U10_Z_31) );
  AND2_X1 U940 ( .A1(in2[1]), .A2(n1563), .ZN(U10_Z_30) );
  AND2_X1 U941 ( .A1(in2[0]), .A2(n1563), .ZN(U10_Z_29) );
  DFF_X2 ops_out_reg_0_ ( .D(U9_Z_0), .CK(clock), .Q(ops_out[0]) );
  DFF_X2 ops_out_reg_1_ ( .D(U9_Z_1), .CK(clock), .Q(ops_out[1]) );
  DFF_X2 ops_out_reg_3_ ( .D(U9_Z_3), .CK(clock), .Q(ops_out[3]) );
  DFF_X2 ops_out_reg_10_ ( .D(U9_Z_10), .CK(clock), .Q(ops_out[10]) );
  DFF_X2 ops_out_reg_11_ ( .D(U9_Z_11), .CK(clock), .Q(ops_out[11]) );
  DFF_X2 ops_out_reg_12_ ( .D(U9_Z_12), .CK(clock), .Q(ops_out[12]) );
  DFF_X2 ops_out_reg_13_ ( .D(U9_Z_13), .CK(clock), .Q(ops_out[13]) );
  DFF_X2 ops_out_reg_14_ ( .D(U9_Z_14), .CK(clock), .Q(ops_out[14]) );
  DFF_X2 ops_out_reg_15_ ( .D(U9_Z_15), .CK(clock), .Q(ops_out[15]) );
  DFF_X2 ops_out_reg_16_ ( .D(U9_Z_16), .CK(clock), .Q(ops_out[16]) );
  DFF_X2 ops_out_reg_17_ ( .D(U9_Z_17), .CK(clock), .Q(ops_out[17]) );
  DFF_X2 ops_out_reg_18_ ( .D(U9_Z_18), .CK(clock), .Q(ops_out[18]) );
  DFF_X2 ops_out_reg_19_ ( .D(U9_Z_19), .CK(clock), .Q(ops_out[19]) );
  DFF_X2 ops_out_reg_20_ ( .D(U9_Z_20), .CK(clock), .Q(ops_out[20]) );
  DFF_X2 ops_out_reg_21_ ( .D(U9_Z_21), .CK(clock), .Q(ops_out[21]) );
  DFF_X2 ops_out_reg_22_ ( .D(U9_Z_22), .CK(clock), .Q(ops_out[22]) );
  DFF_X2 ops_out_reg_23_ ( .D(U9_Z_23), .CK(clock), .Q(ops_out[23]) );
  DFF_X2 ops_out_reg_24_ ( .D(U9_Z_24), .CK(clock), .Q(ops_out[24]) );
  DFF_X2 ops_out_reg_25_ ( .D(U9_Z_25), .CK(clock), .Q(ops_out[25]) );
  DFF_X2 ops_out_reg_26_ ( .D(U9_Z_26), .CK(clock), .Q(ops_out[26]) );
  DFF_X2 ops_out_reg_27_ ( .D(U9_Z_27), .CK(clock), .Q(ops_out[27]) );
  DFF_X2 ops_out_reg_28_ ( .D(U9_Z_28), .CK(clock), .Q(ops_out[28]) );
  DFF_X2 ops_out_reg_29_ ( .D(U9_Z_29), .CK(clock), .Q(ops_out[29]) );
  DFF_X2 ops_out_reg_30_ ( .D(U9_Z_30), .CK(clock), .Q(ops_out[30]) );
  DFF_X2 ops_out_reg_31_ ( .D(U9_Z_31), .CK(clock), .Q(ops_out[31]) );
  DFF_X2 ops_out_reg_8_ ( .D(U9_Z_8), .CK(clock), .Q(ops_out[8]) );
  DFF_X2 ops_out_reg_9_ ( .D(U9_Z_9), .CK(clock), .Q(ops_out[9]) );
  DFF_X2 ops_out_reg_4_ ( .D(U9_Z_4), .CK(clock), .Q(ops_out[4]) );
  DFF_X2 ops_out_reg_5_ ( .D(U9_Z_5), .CK(clock), .Q(ops_out[5]) );
  DFF_X2 ops_out_reg_6_ ( .D(U9_Z_6), .CK(clock), .Q(ops_out[6]) );
  DFF_X2 ops_out_reg_7_ ( .D(U9_Z_7), .CK(clock), .Q(ops_out[7]) );
  DFF_X2 ops_out_reg_2_ ( .D(U9_Z_2), .CK(clock), .Q(ops_out[2]) );
  NOR2_X2 U942 ( .A1(n1494), .A2(n1495), .ZN(n1049) );
  OAI22_X2 U943 ( .A1(n1252), .A2(n1255), .B1(n1496), .B2(n1497), .ZN(n828) );
  OAI22_X2 U944 ( .A1(n1073), .A2(n1076), .B1(n1498), .B2(n1499), .ZN(n787) );
  NAND2_X2 U945 ( .A1(n1500), .A2(n1501), .ZN(n1029) );
  NAND2_X2 U946 ( .A1(n1502), .A2(n1503), .ZN(n1387) );
  NAND2_X2 U947 ( .A1(n1504), .A2(n1505), .ZN(n1208) );
  NAND2_X2 U948 ( .A1(n1506), .A2(n1507), .ZN(n1000) );
  OAI22_X2 U949 ( .A1(n894), .A2(n897), .B1(n1508), .B2(n1509), .ZN(n869) );
  NOR2_X2 U950 ( .A1(n1510), .A2(n1511), .ZN(n1405) );
  NAND2_X2 U951 ( .A1(n1512), .A2(n1513), .ZN(n1365) );
  NOR2_X2 U952 ( .A1(n1514), .A2(n1515), .ZN(n1226) );
  NAND2_X2 U953 ( .A1(n1516), .A2(n1517), .ZN(n1186) );
  NAND2_X2 U954 ( .A1(n1518), .A2(n1519), .ZN(n903) );
  NOR2_X2 U955 ( .A1(n1520), .A2(n1521), .ZN(n932) );
  NAND2_X2 U956 ( .A1(n1522), .A2(n1523), .ZN(n951) );
  NAND2_X2 U957 ( .A1(n1524), .A2(n1525), .ZN(n1275) );
  NOR2_X2 U958 ( .A1(n1526), .A2(n1527), .ZN(n1407) );
  NAND2_X2 U959 ( .A1(n1528), .A2(n1529), .ZN(n1388) );
  NAND2_X2 U960 ( .A1(n1530), .A2(n1531), .ZN(n1358) );
  NAND2_X2 U961 ( .A1(n1532), .A2(n1533), .ZN(n1096) );
  NOR2_X2 U962 ( .A1(n1534), .A2(n1535), .ZN(n1228) );
  NAND2_X2 U963 ( .A1(n1536), .A2(n1537), .ZN(n1209) );
  NAND2_X2 U964 ( .A1(n1538), .A2(n1539), .ZN(n1179) );
  AOI21_X2 U965 ( .B1(U6_B_22_), .B2(U6_A_22_), .A(n973), .ZN(n984) );
  AOI222_X1 U966 ( .A1(n1001), .A2(n992), .B1(U6_B_18_), .B2(U6_A_18_), .C1(
        n859), .C2(n1000), .ZN(n1005) );
  NAND2_X2 U967 ( .A1(n1540), .A2(n1541), .ZN(n917) );
  NAND2_X2 U968 ( .A1(n1542), .A2(n1543), .ZN(n1007) );
  NAND2_X2 U969 ( .A1(n1544), .A2(n1545), .ZN(n1030) );
  NOR2_X2 U970 ( .A1(n1546), .A2(n1547), .ZN(n1047) );
  NAND2_X2 U971 ( .A1(n1548), .A2(n1549), .ZN(n1261) );
  NAND2_X2 U972 ( .A1(n1550), .A2(n1551), .ZN(n1309) );
  NOR2_X2 U973 ( .A1(n1552), .A2(n1553), .ZN(n1290) );
  NAND2_X2 U974 ( .A1(n1554), .A2(n1555), .ZN(n1082) );
  NAND2_X2 U975 ( .A1(n1556), .A2(n1557), .ZN(n1130) );
  NOR2_X2 U976 ( .A1(n1558), .A2(n1559), .ZN(n1111) );
  AOI222_X1 U977 ( .A1(n1359), .A2(n1350), .B1(U5_B_18_), .B2(U5_A_18_), .C1(
        n818), .C2(n1358), .ZN(n1363) );
  AOI21_X2 U978 ( .B1(U5_B_22_), .B2(U5_A_22_), .A(n1331), .ZN(n1342) );
  AOI222_X1 U979 ( .A1(n1180), .A2(n1171), .B1(U4_B_18_), .B2(U4_A_18_), .C1(
        n777), .C2(n1179), .ZN(n1184) );
  AOI21_X2 U980 ( .B1(U4_B_22_), .B2(U4_A_22_), .A(n1152), .ZN(n1163) );
  XOR2_X2 U981 ( .A(in2[18]), .B(in2[14]), .Z(n1487) );
  XOR2_X2 U982 ( .A(in2[19]), .B(in2[15]), .Z(n1485) );
  XOR2_X2 U983 ( .A(in1[20]), .B(in1[29]), .Z(n1450) );
  XOR2_X2 U984 ( .A(in1[21]), .B(in1[30]), .Z(n1448) );
  XOR2_X2 U985 ( .A(in1[22]), .B(in1[31]), .Z(n1446) );
  INV_X4 U986 ( .A(n1563), .ZN(n1560) );
  INV_X4 U987 ( .A(reset), .ZN(n1563) );
  INV_X4 U988 ( .A(n1563), .ZN(n1561) );
  INV_X4 U989 ( .A(n1563), .ZN(n1562) );
  AOI21_X2 U990 ( .B1(n992), .B2(n993), .A(n994), .ZN(n976) );
  AOI21_X2 U991 ( .B1(n1350), .B2(n1351), .A(n1352), .ZN(n1334) );
  AOI21_X2 U992 ( .B1(n1171), .B2(n1172), .A(n1173), .ZN(n1155) );
  OAI21_X2 U993 ( .B1(n1061), .B2(n873), .A(n903), .ZN(n1060) );
  AOI21_X2 U994 ( .B1(n911), .B2(n1062), .A(n908), .ZN(n1061) );
  OAI21_X2 U995 ( .B1(n1419), .B2(n832), .A(n1261), .ZN(n1418) );
  AOI21_X2 U996 ( .B1(n1269), .B2(n1420), .A(n1266), .ZN(n1419) );
  OAI21_X2 U997 ( .B1(n1240), .B2(n791), .A(n1082), .ZN(n1239) );
  AOI21_X2 U998 ( .B1(n1090), .B2(n1241), .A(n1087), .ZN(n1240) );
  OAI21_X2 U999 ( .B1(n953), .B2(n962), .A(n952), .ZN(n959) );
  OAI21_X2 U1000 ( .B1(n1311), .B2(n1320), .A(n1310), .ZN(n1317) );
  OAI21_X2 U1001 ( .B1(n1132), .B2(n1141), .A(n1131), .ZN(n1138) );
  OAI21_X2 U1002 ( .B1(n1025), .B2(n1026), .A(n1027), .ZN(n1024) );
  OAI21_X2 U1003 ( .B1(n1383), .B2(n1384), .A(n1385), .ZN(n1382) );
  OAI21_X2 U1004 ( .B1(n1204), .B2(n1205), .A(n1206), .ZN(n1203) );
  AOI21_X2 U1005 ( .B1(n1058), .B2(n893), .A(n869), .ZN(n1056) );
  AOI21_X2 U1006 ( .B1(n1416), .B2(n1251), .A(n828), .ZN(n1414) );
  AOI21_X2 U1007 ( .B1(n1237), .B2(n1072), .A(n787), .ZN(n1235) );
  OAI21_X2 U1008 ( .B1(n976), .B2(n985), .A(n977), .ZN(n982) );
  OAI21_X2 U1009 ( .B1(n1334), .B2(n1343), .A(n1335), .ZN(n1340) );
  OAI21_X2 U1010 ( .B1(n1155), .B2(n1164), .A(n1156), .ZN(n1161) );
  OAI21_X2 U1011 ( .B1(n939), .B2(n940), .A(n941), .ZN(n936) );
  OAI21_X2 U1012 ( .B1(n1297), .B2(n1298), .A(n1299), .ZN(n1294) );
  OAI21_X2 U1013 ( .B1(n1118), .B2(n1119), .A(n1120), .ZN(n1115) );
  OAI21_X2 U1014 ( .B1(n909), .B2(n910), .A(n911), .ZN(n904) );
  OAI21_X2 U1015 ( .B1(n1267), .B2(n1268), .A(n1269), .ZN(n1262) );
  OAI21_X2 U1016 ( .B1(n1088), .B2(n1089), .A(n1090), .ZN(n1083) );
  AOI21_X2 U1017 ( .B1(n874), .B2(n904), .A(n873), .ZN(n900) );
  AOI21_X2 U1018 ( .B1(n833), .B2(n1262), .A(n832), .ZN(n1258) );
  AOI21_X2 U1019 ( .B1(n792), .B2(n1083), .A(n791), .ZN(n1079) );
  OAI21_X2 U1020 ( .B1(n973), .B2(n977), .A(n978), .ZN(n970) );
  OAI21_X2 U1021 ( .B1(n1331), .B2(n1335), .A(n1336), .ZN(n1328) );
  OAI21_X2 U1022 ( .B1(n1152), .B2(n1156), .A(n1157), .ZN(n1149) );
  OAI211_X2 U1023 ( .C1(n1019), .C2(n1020), .A(n1021), .B(n1022), .ZN(n992) );
  AOI22_X2 U1024 ( .A1(U6_B_15_), .A2(n1023), .B1(U6_A_15_), .B2(n1024), .ZN(
        n1022) );
  OAI211_X2 U1025 ( .C1(n1377), .C2(n1378), .A(n1379), .B(n1380), .ZN(n1350)
         );
  AOI22_X2 U1026 ( .A1(U5_B_15_), .A2(n1381), .B1(U5_A_15_), .B2(n1382), .ZN(
        n1380) );
  OAI211_X2 U1027 ( .C1(n1198), .C2(n1199), .A(n1200), .B(n1201), .ZN(n1171)
         );
  AOI22_X2 U1028 ( .A1(U4_B_15_), .A2(n1202), .B1(U4_A_15_), .B2(n1203), .ZN(
        n1201) );
  AOI22_X2 U1029 ( .A1(U6_A_5_), .A2(U6_B_5_), .B1(n875), .B2(n876), .ZN(n911)
         );
  AOI22_X2 U1030 ( .A1(U5_A_5_), .A2(U5_B_5_), .B1(n834), .B2(n835), .ZN(n1269) );
  AOI22_X2 U1031 ( .A1(U4_A_5_), .A2(U4_B_5_), .B1(n793), .B2(n794), .ZN(n1090) );
  AOI22_X2 U1032 ( .A1(U6_A_13_), .A2(U6_B_13_), .B1(n865), .B2(n866), .ZN(
        n1026) );
  AOI22_X2 U1033 ( .A1(U5_A_13_), .A2(U5_B_13_), .B1(n824), .B2(n825), .ZN(
        n1384) );
  AOI22_X2 U1034 ( .A1(U4_A_13_), .A2(U4_B_13_), .B1(n783), .B2(n784), .ZN(
        n1205) );
  AOI21_X2 U1035 ( .B1(n1065), .B2(U6_A_1_), .A(n879), .ZN(n939) );
  OAI21_X2 U1036 ( .B1(n1065), .B2(U6_A_1_), .A(U6_B_1_), .ZN(n1066) );
  AOI21_X2 U1037 ( .B1(n1423), .B2(U5_A_1_), .A(n838), .ZN(n1297) );
  OAI21_X2 U1038 ( .B1(n1423), .B2(U5_A_1_), .A(U5_B_1_), .ZN(n1424) );
  AOI21_X2 U1039 ( .B1(n1244), .B2(U4_A_1_), .A(n797), .ZN(n1118) );
  OAI21_X2 U1040 ( .B1(n1244), .B2(U4_A_1_), .A(U4_B_1_), .ZN(n1245) );
  OAI211_X2 U1041 ( .C1(n1063), .C2(n941), .A(n938), .B(n1064), .ZN(n916) );
  OAI211_X2 U1042 ( .C1(U6_B_2_), .C2(U6_A_2_), .A(n878), .B(n877), .ZN(n1064)
         );
  OAI211_X2 U1043 ( .C1(n1421), .C2(n1299), .A(n1296), .B(n1422), .ZN(n1274)
         );
  OAI211_X2 U1044 ( .C1(U5_B_2_), .C2(U5_A_2_), .A(n837), .B(n836), .ZN(n1422)
         );
  OAI211_X2 U1045 ( .C1(n1242), .C2(n1120), .A(n1117), .B(n1243), .ZN(n1095)
         );
  OAI211_X2 U1046 ( .C1(U4_B_2_), .C2(U4_A_2_), .A(n796), .B(n795), .ZN(n1243)
         );
  AOI21_X2 U1047 ( .B1(n931), .B2(n926), .A(n844), .ZN(n929) );
  AOI21_X2 U1048 ( .B1(n1110), .B2(n1105), .A(n762), .ZN(n1108) );
  OAI21_X2 U1049 ( .B1(U6_A_23_), .B2(U6_B_23_), .A(n856), .ZN(n975) );
  OAI21_X2 U1050 ( .B1(U5_A_23_), .B2(U5_B_23_), .A(n815), .ZN(n1333) );
  OAI21_X2 U1051 ( .B1(U4_A_23_), .B2(U4_B_23_), .A(n774), .ZN(n1154) );
  AOI21_X2 U1052 ( .B1(n1289), .B2(n1284), .A(n803), .ZN(n1287) );
  AOI21_X2 U1053 ( .B1(n959), .B2(n951), .A(n848), .ZN(n957) );
  AOI21_X2 U1054 ( .B1(U6_B_29_), .B2(U6_A_29_), .A(n933), .ZN(n943) );
  AOI21_X2 U1055 ( .B1(n926), .B2(n846), .A(n932), .ZN(n944) );
  AOI21_X2 U1056 ( .B1(n1317), .B2(n1309), .A(n807), .ZN(n1315) );
  AOI21_X2 U1057 ( .B1(U5_B_29_), .B2(U5_A_29_), .A(n1291), .ZN(n1301) );
  AOI21_X2 U1058 ( .B1(n1284), .B2(n805), .A(n1290), .ZN(n1302) );
  AOI21_X2 U1059 ( .B1(n1138), .B2(n1130), .A(n766), .ZN(n1136) );
  AOI21_X2 U1060 ( .B1(U4_B_29_), .B2(U4_A_29_), .A(n1112), .ZN(n1122) );
  AOI21_X2 U1061 ( .B1(n1105), .B2(n764), .A(n1111), .ZN(n1123) );
  AOI22_X2 U1062 ( .A1(U4_A_21_), .A2(U4_B_21_), .B1(n772), .B2(n773), .ZN(
        n1156) );
  AOI22_X2 U1063 ( .A1(U6_A_17_), .A2(U6_B_17_), .B1(n860), .B2(n861), .ZN(
        n997) );
  AOI22_X2 U1064 ( .A1(U5_A_17_), .A2(U5_B_17_), .B1(n819), .B2(n820), .ZN(
        n1355) );
  AOI22_X2 U1065 ( .A1(U4_A_17_), .A2(U4_B_17_), .B1(n778), .B2(n779), .ZN(
        n1176) );
  AOI21_X2 U1066 ( .B1(U6_A_25_), .B2(U6_B_25_), .A(n955), .ZN(n964) );
  OAI21_X2 U1067 ( .B1(n954), .B2(n953), .A(n966), .ZN(n965) );
  AOI21_X2 U1068 ( .B1(U5_A_25_), .B2(U5_B_25_), .A(n1313), .ZN(n1322) );
  OAI21_X2 U1069 ( .B1(n1312), .B2(n1311), .A(n1324), .ZN(n1323) );
  AOI21_X2 U1070 ( .B1(U4_A_25_), .B2(U4_B_25_), .A(n1134), .ZN(n1143) );
  OAI21_X2 U1071 ( .B1(n1133), .B2(n1132), .A(n1145), .ZN(n1144) );
  AOI22_X2 U1072 ( .A1(U6_A_21_), .A2(U6_B_21_), .B1(n854), .B2(n855), .ZN(
        n977) );
  AOI22_X2 U1073 ( .A1(U5_A_21_), .A2(U5_B_21_), .B1(n813), .B2(n814), .ZN(
        n1335) );
  AOI21_X2 U1074 ( .B1(n1034), .B2(n863), .A(n864), .ZN(n1032) );
  AOI21_X2 U1075 ( .B1(n1392), .B2(n822), .A(n823), .ZN(n1390) );
  AOI21_X2 U1076 ( .B1(n1213), .B2(n781), .A(n782), .ZN(n1211) );
  OAI21_X2 U1077 ( .B1(n853), .B2(n973), .A(n978), .ZN(n980) );
  OAI21_X2 U1078 ( .B1(n812), .B2(n1331), .A(n1336), .ZN(n1338) );
  OAI21_X2 U1079 ( .B1(n771), .B2(n1152), .A(n1157), .ZN(n1159) );
  AOI21_X2 U1080 ( .B1(U6_B_13_), .B2(U6_A_13_), .A(n1039), .ZN(n1041) );
  AOI21_X2 U1081 ( .B1(n1038), .B2(n1030), .A(n866), .ZN(n1042) );
  AOI21_X2 U1082 ( .B1(U6_B_17_), .B2(U6_A_17_), .A(n1012), .ZN(n1014) );
  AOI21_X2 U1083 ( .B1(n1007), .B2(n992), .A(n861), .ZN(n1015) );
  AOI21_X2 U1084 ( .B1(U6_B_9_), .B2(U6_A_9_), .A(n894), .ZN(n891) );
  AOI21_X2 U1085 ( .B1(n893), .B2(n872), .A(n871), .ZN(n892) );
  AOI21_X2 U1086 ( .B1(U5_B_9_), .B2(U5_A_9_), .A(n1252), .ZN(n1249) );
  AOI21_X2 U1087 ( .B1(n1251), .B2(n831), .A(n830), .ZN(n1250) );
  AOI21_X2 U1088 ( .B1(U5_B_13_), .B2(U5_A_13_), .A(n1397), .ZN(n1399) );
  AOI21_X2 U1089 ( .B1(n1396), .B2(n1388), .A(n825), .ZN(n1400) );
  AOI21_X2 U1090 ( .B1(U5_B_17_), .B2(U5_A_17_), .A(n1370), .ZN(n1372) );
  AOI21_X2 U1091 ( .B1(n1365), .B2(n1350), .A(n820), .ZN(n1373) );
  AOI21_X2 U1092 ( .B1(U4_B_9_), .B2(U4_A_9_), .A(n1073), .ZN(n1070) );
  AOI21_X2 U1093 ( .B1(n1072), .B2(n790), .A(n789), .ZN(n1071) );
  AOI21_X2 U1094 ( .B1(U4_B_13_), .B2(U4_A_13_), .A(n1218), .ZN(n1220) );
  AOI21_X2 U1095 ( .B1(n1217), .B2(n1209), .A(n784), .ZN(n1221) );
  AOI21_X2 U1096 ( .B1(U4_B_17_), .B2(U4_A_17_), .A(n1191), .ZN(n1193) );
  AOI21_X2 U1097 ( .B1(n1186), .B2(n1171), .A(n779), .ZN(n1194) );
  AOI21_X2 U1098 ( .B1(U6_A_21_), .B2(U6_B_21_), .A(n974), .ZN(n987) );
  OAI21_X2 U1099 ( .B1(n972), .B2(n976), .A(n989), .ZN(n988) );
  AOI21_X2 U1100 ( .B1(U5_A_21_), .B2(U5_B_21_), .A(n1332), .ZN(n1345) );
  OAI21_X2 U1101 ( .B1(n1330), .B2(n1334), .A(n1347), .ZN(n1346) );
  AOI21_X2 U1102 ( .B1(U4_A_21_), .B2(U4_B_21_), .A(n1153), .ZN(n1166) );
  OAI21_X2 U1103 ( .B1(n1151), .B2(n1155), .A(n1168), .ZN(n1167) );
  AOI22_X2 U1104 ( .A1(U6_A_25_), .A2(U6_B_25_), .B1(n850), .B2(n851), .ZN(
        n952) );
  AOI22_X2 U1105 ( .A1(U5_A_25_), .A2(U5_B_25_), .B1(n809), .B2(n810), .ZN(
        n1310) );
  AOI22_X2 U1106 ( .A1(U4_A_25_), .A2(U4_B_25_), .B1(n768), .B2(n769), .ZN(
        n1131) );
  AOI22_X2 U1107 ( .A1(U6_A_29_), .A2(U6_B_29_), .B1(n845), .B2(n932), .ZN(
        n924) );
  AOI22_X2 U1108 ( .A1(U5_A_29_), .A2(U5_B_29_), .B1(n804), .B2(n1290), .ZN(
        n1282) );
  AOI22_X2 U1109 ( .A1(U4_A_29_), .A2(U4_B_29_), .B1(n763), .B2(n1111), .ZN(
        n1103) );
  AOI21_X2 U1110 ( .B1(U6_A_5_), .B2(U6_B_5_), .A(n909), .ZN(n913) );
  AOI21_X2 U1111 ( .B1(U5_A_5_), .B2(U5_B_5_), .A(n1267), .ZN(n1271) );
  AOI21_X2 U1112 ( .B1(U4_A_5_), .B2(U4_B_5_), .A(n1088), .ZN(n1092) );
  AOI211_X2 U1113 ( .C1(n842), .C2(n839), .A(n1560), .B(n1423), .ZN(U7_Z_0) );
  AOI211_X2 U1114 ( .C1(n801), .C2(n798), .A(n1562), .B(n1244), .ZN(U8_Z_0) );
  AOI211_X2 U1115 ( .C1(n880), .C2(n883), .A(n1561), .B(n1065), .ZN(U9_Z_0) );
  OAI21_X2 U1116 ( .B1(U6_A_2_), .B2(U6_B_2_), .A(n941), .ZN(n1003) );
  OAI21_X2 U1117 ( .B1(U5_A_2_), .B2(U5_B_2_), .A(n1299), .ZN(n1361) );
  OAI21_X2 U1118 ( .B1(U4_A_2_), .B2(U4_B_2_), .A(n1120), .ZN(n1182) );
endmodule

