
module w_op ( clock, reset, in1, in2, in3, in4, ops_out );
  input [31:0] in1;
  input [31:0] in2;
  input [31:0] in3;
  input [31:0] in4;
  output [31:0] ops_out;
  input clock, reset;
  wire   U7_Z_0, U7_Z_1, U7_Z_2, U7_Z_3, U7_Z_4, U7_Z_5, U7_Z_6, U7_Z_7,
         U7_Z_8, U7_Z_9, U7_Z_10, U7_Z_11, U7_Z_12, U7_Z_13, U7_Z_14, U7_Z_15,
         U7_Z_16, U7_Z_17, U7_Z_18, U7_Z_19, U7_Z_20, U7_Z_21, U7_Z_22,
         U7_Z_23, U7_Z_24, U7_Z_25, U7_Z_26, U7_Z_27, U7_Z_28, U7_Z_29,
         U7_Z_30, U7_Z_31, n366, n368, n370, n371, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n385, n386, n387, n388, n389,
         n390, n392, n393, n394, n395, n396, n397, n398, n400, n401, n402,
         n403, n404, n406, n407, n408, n409, n410, n411, n412, n413, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n488, n489, n491, n492, n493, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111;

  NOR2_X2 U3 ( .A1(n1110), .A2(n506), .ZN(U7_Z_9) );
  XOR2_X2 U4 ( .A(n507), .B(n508), .Z(n506) );
  NOR2_X2 U7 ( .A1(n1110), .A2(n515), .ZN(U7_Z_8) );
  XOR2_X2 U8 ( .A(n509), .B(n516), .Z(n515) );
  NOR2_X2 U10 ( .A1(n1110), .A2(n517), .ZN(U7_Z_7) );
  XNOR2_X2 U11 ( .A(n518), .B(n519), .ZN(n517) );
  NAND2_X2 U12 ( .A1(n520), .A2(n521), .ZN(n519) );
  NOR2_X2 U14 ( .A1(n1110), .A2(n525), .ZN(U7_Z_6) );
  XOR2_X2 U15 ( .A(n522), .B(n526), .Z(n525) );
  NOR2_X2 U17 ( .A1(n1110), .A2(n528), .ZN(U7_Z_5) );
  XOR2_X2 U18 ( .A(n529), .B(n530), .Z(n528) );
  NAND2_X2 U19 ( .A1(n531), .A2(n527), .ZN(n530) );
  NAND2_X2 U20 ( .A1(n532), .A2(n533), .ZN(n527) );
  NOR2_X2 U22 ( .A1(n1110), .A2(n537), .ZN(U7_Z_4) );
  XOR2_X2 U23 ( .A(n532), .B(n538), .Z(n537) );
  NAND2_X2 U24 ( .A1(n531), .A2(n533), .ZN(n538) );
  NOR2_X2 U25 ( .A1(n1110), .A2(n539), .ZN(U7_Z_31) );
  XOR2_X2 U26 ( .A(n540), .B(n541), .Z(n539) );
  XOR2_X2 U27 ( .A(n542), .B(n543), .Z(n541) );
  XOR2_X2 U28 ( .A(n544), .B(n545), .Z(n543) );
  NOR3_X2 U30 ( .A1(n547), .A2(n548), .A3(n549), .ZN(n546) );
  OAI221_X2 U33 ( .B1(n553), .B2(n497), .C1(n554), .C2(n434), .A(n555), .ZN(
        n544) );
  NAND4_X2 U34 ( .A1(n556), .A2(n557), .A3(n558), .A4(n437), .ZN(n555) );
  NAND2_X2 U35 ( .A1(n434), .A2(n497), .ZN(n557) );
  NOR2_X2 U36 ( .A1(in1[8]), .A2(n435), .ZN(n553) );
  NAND4_X2 U39 ( .A1(n564), .A2(n565), .A3(n374), .A4(n566), .ZN(n561) );
  NAND2_X2 U40 ( .A1(n563), .A2(n560), .ZN(n565) );
  XOR2_X2 U41 ( .A(n567), .B(n568), .Z(n540) );
  XNOR2_X2 U42 ( .A(in3[31]), .B(in1[9]), .ZN(n568) );
  XNOR2_X2 U43 ( .A(in4[31]), .B(in2[2]), .ZN(n567) );
  NOR2_X2 U44 ( .A1(n1110), .A2(n569), .ZN(U7_Z_30) );
  XOR2_X2 U45 ( .A(n563), .B(n570), .Z(n569) );
  XNOR2_X2 U46 ( .A(n571), .B(n560), .ZN(n570) );
  XNOR2_X2 U47 ( .A(n572), .B(n573), .ZN(n560) );
  XOR2_X2 U48 ( .A(in4[30]), .B(in2[1]), .Z(n573) );
  NAND2_X2 U49 ( .A1(n552), .A2(n574), .ZN(n572) );
  NAND3_X2 U50 ( .A1(n496), .A2(n447), .A3(n550), .ZN(n574) );
  NAND2_X2 U52 ( .A1(n559), .A2(n576), .ZN(n571) );
  NAND3_X2 U53 ( .A1(n374), .A2(n566), .A3(n564), .ZN(n576) );
  XNOR2_X2 U55 ( .A(n581), .B(n582), .ZN(n563) );
  XOR2_X2 U58 ( .A(n497), .B(in1[8]), .Z(n581) );
  NOR2_X2 U59 ( .A1(n1110), .A2(n585), .ZN(U7_Z_3) );
  XOR2_X2 U60 ( .A(n586), .B(n587), .Z(n585) );
  NAND2_X2 U61 ( .A1(n427), .A2(n588), .ZN(n587) );
  NOR2_X2 U63 ( .A1(n592), .A2(n593), .ZN(n590) );
  NOR2_X2 U64 ( .A1(n1110), .A2(n594), .ZN(U7_Z_29) );
  XOR2_X2 U65 ( .A(n595), .B(n596), .Z(n594) );
  NOR2_X2 U68 ( .A1(n577), .A2(n578), .ZN(n580) );
  XOR2_X2 U69 ( .A(n597), .B(n598), .Z(n577) );
  NAND2_X2 U72 ( .A1(n498), .A2(n436), .ZN(n558) );
  XNOR2_X2 U73 ( .A(n600), .B(n601), .ZN(n578) );
  NOR2_X2 U76 ( .A1(in4[29]), .A2(in2[0]), .ZN(n549) );
  NOR2_X2 U77 ( .A1(n1110), .A2(n602), .ZN(U7_Z_28) );
  XOR2_X2 U78 ( .A(n564), .B(n603), .Z(n602) );
  NOR2_X2 U80 ( .A1(n604), .A2(n605), .ZN(n579) );
  NAND2_X2 U81 ( .A1(n605), .A2(n604), .ZN(n566) );
  XNOR2_X2 U82 ( .A(n550), .B(n606), .ZN(n604) );
  NOR2_X2 U83 ( .A1(n575), .A2(n548), .ZN(n606) );
  NOR2_X2 U84 ( .A1(in2[31]), .A2(in4[28]), .ZN(n548) );
  OAI221_X2 U86 ( .B1(in4[27]), .B2(in2[30]), .C1(n610), .C2(n451), .A(n464), 
        .ZN(n609) );
  NOR3_X2 U87 ( .A1(n456), .A2(n612), .A3(n613), .ZN(n610) );
  XNOR2_X2 U89 ( .A(n556), .B(n614), .ZN(n605) );
  NOR2_X2 U90 ( .A1(n584), .A2(n599), .ZN(n614) );
  NOR2_X2 U91 ( .A1(in1[6]), .A2(in3[28]), .ZN(n599) );
  OAI221_X2 U93 ( .B1(in3[27]), .B2(in1[5]), .C1(n618), .C2(n441), .A(n439), 
        .ZN(n617) );
  NOR3_X2 U94 ( .A1(n375), .A2(n620), .A3(n621), .ZN(n618) );
  OAI221_X2 U97 ( .B1(n624), .B2(n625), .C1(n626), .C2(n627), .A(n628), .ZN(
        n623) );
  NOR3_X2 U98 ( .A1(n629), .A2(n630), .A3(n376), .ZN(n626) );
  NOR2_X2 U100 ( .A1(n1110), .A2(n632), .ZN(U7_Z_27) );
  XNOR2_X2 U101 ( .A(n625), .B(n633), .ZN(n632) );
  XOR2_X2 U102 ( .A(n634), .B(n450), .Z(n633) );
  XOR2_X2 U103 ( .A(n635), .B(n636), .Z(n624) );
  XOR2_X2 U105 ( .A(in4[27]), .B(n463), .Z(n635) );
  XOR2_X2 U107 ( .A(n640), .B(n641), .Z(n625) );
  XOR2_X2 U109 ( .A(in3[27]), .B(n438), .Z(n640) );
  NOR2_X2 U110 ( .A1(n1110), .A2(n644), .ZN(U7_Z_26) );
  XOR2_X2 U111 ( .A(n639), .B(n645), .Z(n644) );
  NAND2_X2 U112 ( .A1(n628), .A2(n371), .ZN(n645) );
  NOR2_X2 U113 ( .A1(n646), .A2(n647), .ZN(n631) );
  NAND2_X2 U114 ( .A1(n647), .A2(n646), .ZN(n628) );
  XNOR2_X2 U115 ( .A(n642), .B(n648), .ZN(n646) );
  NOR2_X2 U116 ( .A1(n440), .A2(n643), .ZN(n648) );
  NOR2_X2 U117 ( .A1(in1[4]), .A2(in3[26]), .ZN(n643) );
  NAND2_X2 U118 ( .A1(in3[26]), .A2(in1[4]), .ZN(n615) );
  NAND2_X2 U121 ( .A1(n442), .A2(n443), .ZN(n649) );
  XNOR2_X2 U122 ( .A(n637), .B(n650), .ZN(n647) );
  NOR2_X2 U123 ( .A1(n465), .A2(n638), .ZN(n650) );
  NOR2_X2 U124 ( .A1(in2[29]), .A2(in4[26]), .ZN(n638) );
  NAND2_X2 U125 ( .A1(in4[26]), .A2(in2[29]), .ZN(n607) );
  NAND2_X2 U128 ( .A1(n468), .A2(n453), .ZN(n651) );
  OAI22_X2 U130 ( .A1(n654), .A2(n655), .B1(n376), .B2(n656), .ZN(n627) );
  NOR2_X2 U131 ( .A1(n1110), .A2(n658), .ZN(U7_Z_25) );
  XOR2_X2 U132 ( .A(n659), .B(n660), .Z(n658) );
  NAND2_X2 U135 ( .A1(n654), .A2(n655), .ZN(n657) );
  XNOR2_X2 U136 ( .A(n661), .B(n662), .ZN(n655) );
  NOR2_X2 U138 ( .A1(in4[25]), .A2(in2[28]), .ZN(n613) );
  XOR2_X2 U140 ( .A(n663), .B(n664), .Z(n654) );
  NOR2_X2 U143 ( .A1(in3[25]), .A2(in1[3]), .ZN(n621) );
  NOR2_X2 U144 ( .A1(n1110), .A2(n667), .ZN(U7_Z_24) );
  XOR2_X2 U145 ( .A(n629), .B(n668), .Z(n667) );
  NAND2_X2 U147 ( .A1(n669), .A2(n670), .ZN(n656) );
  NOR2_X2 U148 ( .A1(n670), .A2(n669), .ZN(n630) );
  XOR2_X2 U149 ( .A(n671), .B(n456), .Z(n669) );
  OAI221_X2 U150 ( .B1(n461), .B2(n673), .C1(n674), .C2(n503), .A(n675), .ZN(
        n672) );
  NAND4_X2 U151 ( .A1(n473), .A2(n466), .A3(n470), .A4(n676), .ZN(n675) );
  NOR2_X2 U152 ( .A1(n461), .A2(n677), .ZN(n676) );
  NAND2_X2 U154 ( .A1(n652), .A2(n453), .ZN(n671) );
  NOR2_X2 U155 ( .A1(n681), .A2(in4[24]), .ZN(n612) );
  NAND2_X2 U156 ( .A1(in4[24]), .A2(n681), .ZN(n652) );
  XOR2_X2 U157 ( .A(in2[27]), .B(in2[31]), .Z(n681) );
  XOR2_X2 U158 ( .A(n682), .B(n375), .Z(n670) );
  OAI221_X2 U159 ( .B1(n683), .B2(n684), .C1(n445), .C2(n499), .A(n685), .ZN(
        n665) );
  NAND4_X2 U160 ( .A1(n396), .A2(n686), .A3(n380), .A4(n687), .ZN(n685) );
  NOR2_X2 U161 ( .A1(n683), .A2(n688), .ZN(n687) );
  NAND2_X2 U163 ( .A1(n666), .A2(n443), .ZN(n682) );
  NOR2_X2 U164 ( .A1(in1[2]), .A2(in3[24]), .ZN(n620) );
  NAND2_X2 U165 ( .A1(in3[24]), .A2(in1[2]), .ZN(n666) );
  AOI221_X2 U166 ( .B1(n690), .B2(n691), .C1(n366), .C2(n692), .A(n693), .ZN(
        n629) );
  AND4_X2 U167 ( .A1(n694), .A2(n695), .A3(n696), .A4(n697), .ZN(n693) );
  NAND2_X2 U169 ( .A1(n455), .A2(n699), .ZN(n690) );
  NOR2_X2 U171 ( .A1(n1110), .A2(n702), .ZN(U7_Z_23) );
  XOR2_X2 U172 ( .A(n691), .B(n703), .Z(n702) );
  XOR2_X2 U173 ( .A(n692), .B(n704), .Z(n703) );
  XOR2_X2 U175 ( .A(n706), .B(n707), .Z(n692) );
  NAND2_X2 U178 ( .A1(n674), .A2(n503), .ZN(n680) );
  XOR2_X2 U179 ( .A(n476), .B(in2[30]), .Z(n674) );
  XNOR2_X2 U180 ( .A(n710), .B(n711), .ZN(n691) );
  NOR2_X2 U183 ( .A1(in3[23]), .A2(in1[1]), .ZN(n683) );
  NOR2_X2 U184 ( .A1(n1110), .A2(n714), .ZN(U7_Z_22) );
  XOR2_X2 U185 ( .A(n705), .B(n715), .Z(n714) );
  NOR2_X2 U187 ( .A1(n716), .A2(n717), .ZN(n701) );
  NAND2_X2 U188 ( .A1(n717), .A2(n716), .ZN(n695) );
  XOR2_X2 U189 ( .A(n718), .B(n712), .Z(n716) );
  NAND2_X2 U192 ( .A1(n380), .A2(n396), .ZN(n719) );
  NAND2_X2 U193 ( .A1(n686), .A2(n713), .ZN(n718) );
  NAND2_X2 U194 ( .A1(in3[22]), .A2(in1[0]), .ZN(n713) );
  XNOR2_X2 U195 ( .A(n708), .B(n722), .ZN(n717) );
  NOR2_X2 U196 ( .A1(n678), .A2(n709), .ZN(n722) );
  NOR2_X2 U197 ( .A1(n723), .A2(in4[22]), .ZN(n709) );
  XOR2_X2 U198 ( .A(in2[25]), .B(in2[29]), .Z(n723) );
  NAND2_X2 U201 ( .A1(n470), .A2(n473), .ZN(n724) );
  OAI22_X2 U203 ( .A1(n729), .A2(n730), .B1(n379), .B2(n389), .ZN(n700) );
  NAND2_X2 U204 ( .A1(n696), .A2(n694), .ZN(n728) );
  NOR2_X2 U205 ( .A1(n1110), .A2(n731), .ZN(U7_Z_21) );
  XOR2_X2 U206 ( .A(n732), .B(n733), .Z(n731) );
  NAND2_X2 U209 ( .A1(n729), .A2(n730), .ZN(n696) );
  XNOR2_X2 U210 ( .A(n735), .B(n736), .ZN(n730) );
  NOR2_X2 U212 ( .A1(n725), .A2(in4[21]), .ZN(n727) );
  XOR2_X2 U213 ( .A(in2[24]), .B(in2[28]), .Z(n725) );
  XNOR2_X2 U215 ( .A(n738), .B(n739), .ZN(n729) );
  NOR2_X2 U217 ( .A1(in3[21]), .A2(in1[31]), .ZN(n721) );
  NOR2_X2 U219 ( .A1(n1110), .A2(n741), .ZN(U7_Z_20) );
  XOR2_X2 U220 ( .A(n698), .B(n742), .Z(n741) );
  NOR2_X2 U221 ( .A1(n388), .A2(n734), .ZN(n742) );
  NOR2_X2 U222 ( .A1(n743), .A2(n744), .ZN(n734) );
  NAND2_X2 U223 ( .A1(n744), .A2(n743), .ZN(n694) );
  XNOR2_X2 U224 ( .A(n745), .B(n677), .ZN(n743) );
  OAI221_X2 U226 ( .B1(n748), .B2(n749), .C1(n481), .C2(n750), .A(n751), .ZN(
        n747) );
  NAND2_X2 U227 ( .A1(n479), .A2(n475), .ZN(n750) );
  NAND2_X2 U228 ( .A1(n726), .A2(n473), .ZN(n745) );
  NOR2_X2 U229 ( .A1(n753), .A2(in4[20]), .ZN(n737) );
  NAND2_X2 U230 ( .A1(in4[20]), .A2(n753), .ZN(n726) );
  XOR2_X2 U231 ( .A(in2[23]), .B(in2[27]), .Z(n753) );
  XNOR2_X2 U232 ( .A(n754), .B(n688), .ZN(n744) );
  OAI221_X2 U234 ( .B1(n758), .B2(n759), .C1(n760), .C2(n761), .A(n762), .ZN(
        n757) );
  NAND2_X2 U235 ( .A1(n407), .A2(n403), .ZN(n761) );
  NAND2_X2 U236 ( .A1(n720), .A2(n396), .ZN(n754) );
  NOR2_X2 U237 ( .A1(in1[30]), .A2(in3[20]), .ZN(n740) );
  NAND2_X2 U238 ( .A1(in3[20]), .A2(in1[30]), .ZN(n720) );
  OAI221_X2 U240 ( .B1(n767), .B2(n768), .C1(n769), .C2(n770), .A(n771), .ZN(
        n766) );
  NAND2_X2 U241 ( .A1(n386), .A2(n387), .ZN(n770) );
  NOR2_X2 U242 ( .A1(n772), .A2(n767), .ZN(n765) );
  NOR2_X2 U243 ( .A1(n1110), .A2(n773), .ZN(U7_Z_2) );
  XOR2_X2 U244 ( .A(n429), .B(n774), .Z(n773) );
  NOR2_X2 U246 ( .A1(n1110), .A2(n775), .ZN(U7_Z_19) );
  XOR2_X2 U247 ( .A(n776), .B(n777), .Z(n775) );
  NAND2_X2 U248 ( .A1(n387), .A2(n771), .ZN(n777) );
  NAND2_X2 U249 ( .A1(n778), .A2(n779), .ZN(n771) );
  NOR2_X2 U250 ( .A1(n779), .A2(n778), .ZN(n767) );
  XOR2_X2 U251 ( .A(n780), .B(n781), .Z(n778) );
  AOI221_X2 U252 ( .B1(n763), .B2(n755), .C1(n411), .C2(n407), .A(n406), .ZN(
        n781) );
  NOR3_X2 U253 ( .A1(n782), .A2(n783), .A3(n784), .ZN(n763) );
  NAND2_X2 U254 ( .A1(n403), .A2(n762), .ZN(n780) );
  NAND2_X2 U255 ( .A1(in3[19]), .A2(in1[29]), .ZN(n762) );
  NOR2_X2 U256 ( .A1(in1[29]), .A2(in3[19]), .ZN(n758) );
  XOR2_X2 U257 ( .A(n785), .B(n786), .Z(n779) );
  AOI221_X2 U258 ( .B1(n752), .B2(n457), .C1(n787), .C2(n479), .A(n480), .ZN(
        n786) );
  NOR3_X2 U259 ( .A1(n788), .A2(n789), .A3(n482), .ZN(n752) );
  NAND2_X2 U260 ( .A1(n475), .A2(n751), .ZN(n785) );
  NAND2_X2 U261 ( .A1(in4[19]), .A2(n790), .ZN(n751) );
  NOR2_X2 U262 ( .A1(n790), .A2(in4[19]), .ZN(n748) );
  OAI221_X2 U264 ( .B1(n791), .B2(n769), .C1(n381), .C2(n772), .A(n768), .ZN(
        n776) );
  NAND3_X2 U265 ( .A1(n386), .A2(n792), .A3(n385), .ZN(n772) );
  NOR2_X2 U266 ( .A1(n1110), .A2(n793), .ZN(U7_Z_18) );
  XOR2_X2 U267 ( .A(n794), .B(n795), .Z(n793) );
  NAND2_X2 U268 ( .A1(n768), .A2(n386), .ZN(n795) );
  NOR2_X2 U269 ( .A1(n796), .A2(n797), .ZN(n791) );
  NAND2_X2 U270 ( .A1(n797), .A2(n796), .ZN(n768) );
  XOR2_X2 U271 ( .A(n798), .B(n799), .Z(n796) );
  NOR2_X2 U272 ( .A1(n788), .A2(n480), .ZN(n799) );
  NAND2_X2 U273 ( .A1(in4[18]), .A2(n800), .ZN(n749) );
  NOR2_X2 U274 ( .A1(n800), .A2(in4[18]), .ZN(n788) );
  XOR2_X2 U275 ( .A(in2[21]), .B(in2[25]), .Z(n800) );
  NAND2_X2 U276 ( .A1(n481), .A2(n801), .ZN(n798) );
  NAND3_X2 U277 ( .A1(n485), .A2(n457), .A3(n802), .ZN(n801) );
  OAI22_X2 U278 ( .A1(n803), .A2(n504), .B1(n482), .B2(n804), .ZN(n787) );
  XOR2_X2 U279 ( .A(n805), .B(n806), .Z(n797) );
  NOR2_X2 U280 ( .A1(n782), .A2(n406), .ZN(n806) );
  NAND2_X2 U281 ( .A1(in3[18]), .A2(in1[28]), .ZN(n759) );
  NOR2_X2 U282 ( .A1(in1[28]), .A2(in3[18]), .ZN(n782) );
  NAND2_X2 U283 ( .A1(n760), .A2(n807), .ZN(n805) );
  NAND3_X2 U284 ( .A1(n416), .A2(n755), .A3(n412), .ZN(n807) );
  NAND2_X2 U286 ( .A1(n769), .A2(n809), .ZN(n794) );
  NAND3_X2 U287 ( .A1(n792), .A2(n764), .A3(n385), .ZN(n809) );
  NOR2_X2 U289 ( .A1(n1110), .A2(n814), .ZN(U7_Z_17) );
  XOR2_X2 U290 ( .A(n815), .B(n816), .Z(n814) );
  NOR2_X2 U293 ( .A1(n810), .A2(n811), .ZN(n813) );
  XNOR2_X2 U294 ( .A(n817), .B(n818), .ZN(n810) );
  NOR2_X2 U297 ( .A1(in3[17]), .A2(in1[27]), .ZN(n784) );
  XOR2_X2 U298 ( .A(n819), .B(n820), .Z(n811) );
  NAND2_X2 U301 ( .A1(n803), .A2(n504), .ZN(n802) );
  XNOR2_X2 U302 ( .A(in2[20]), .B(in2[24]), .ZN(n803) );
  NOR2_X2 U303 ( .A1(n1110), .A2(n821), .ZN(U7_Z_16) );
  XOR2_X2 U304 ( .A(n764), .B(n822), .Z(n821) );
  NOR2_X2 U306 ( .A1(n823), .A2(n824), .ZN(n812) );
  NAND2_X2 U307 ( .A1(n824), .A2(n823), .ZN(n792) );
  XNOR2_X2 U308 ( .A(n457), .B(n825), .ZN(n823) );
  NOR2_X2 U309 ( .A1(n484), .A2(n789), .ZN(n825) );
  NOR2_X2 U310 ( .A1(n826), .A2(in4[16]), .ZN(n789) );
  NAND2_X2 U311 ( .A1(in4[16]), .A2(n826), .ZN(n804) );
  XOR2_X2 U312 ( .A(in2[19]), .B(in2[23]), .Z(n826) );
  OAI22_X2 U314 ( .A1(n458), .A2(n831), .B1(n460), .B2(n832), .ZN(n830) );
  AND4_X2 U316 ( .A1(n838), .A2(n833), .A3(n839), .A4(n840), .ZN(n829) );
  NOR4_X2 U317 ( .A1(n831), .A2(n841), .A3(n842), .A4(n835), .ZN(n833) );
  XNOR2_X2 U318 ( .A(n755), .B(n843), .ZN(n824) );
  NOR2_X2 U319 ( .A1(n808), .A2(n783), .ZN(n843) );
  NOR2_X2 U320 ( .A1(in1[26]), .A2(in3[16]), .ZN(n783) );
  NAND4_X2 U324 ( .A1(n853), .A2(n848), .A3(n854), .A4(n402), .ZN(n844) );
  AND4_X2 U325 ( .A1(n847), .A2(n855), .A3(n395), .A4(n390), .ZN(n848) );
  NAND2_X2 U328 ( .A1(n862), .A2(n454), .ZN(n860) );
  NAND4_X2 U330 ( .A1(n868), .A2(n869), .A3(n393), .A4(n863), .ZN(n856) );
  NOR2_X2 U332 ( .A1(n1110), .A2(n870), .ZN(U7_Z_15) );
  XOR2_X2 U333 ( .A(n859), .B(n871), .Z(n870) );
  XOR2_X2 U334 ( .A(n861), .B(n872), .Z(n871) );
  XOR2_X2 U336 ( .A(n874), .B(n875), .Z(n861) );
  NOR2_X2 U338 ( .A1(n828), .A2(in4[15]), .ZN(n831) );
  XNOR2_X2 U341 ( .A(n877), .B(n878), .ZN(n859) );
  NAND2_X2 U344 ( .A1(n500), .A2(n420), .ZN(n847) );
  NOR2_X2 U345 ( .A1(n1110), .A2(n880), .ZN(U7_Z_14) );
  XOR2_X2 U346 ( .A(n873), .B(n881), .Z(n880) );
  NOR2_X2 U348 ( .A1(n882), .A2(n883), .ZN(n865) );
  NAND2_X2 U349 ( .A1(n883), .A2(n882), .ZN(n863) );
  XNOR2_X2 U350 ( .A(n884), .B(n879), .ZN(n882) );
  NAND3_X2 U351 ( .A1(n855), .A2(n395), .A3(n886), .ZN(n885) );
  NAND2_X2 U353 ( .A1(n390), .A2(n852), .ZN(n884) );
  NAND2_X2 U354 ( .A1(in3[14]), .A2(n889), .ZN(n852) );
  NOR2_X2 U355 ( .A1(n889), .A2(in3[14]), .ZN(n850) );
  XOR2_X2 U356 ( .A(in1[24]), .B(in1[31]), .Z(n889) );
  XNOR2_X2 U357 ( .A(n890), .B(n876), .ZN(n883) );
  NAND3_X2 U358 ( .A1(n459), .A2(n462), .A3(n892), .ZN(n891) );
  NAND2_X2 U361 ( .A1(in4[14]), .A2(n895), .ZN(n837) );
  NOR2_X2 U362 ( .A1(n895), .A2(in4[14]), .ZN(n835) );
  XOR2_X2 U363 ( .A(in2[17]), .B(in2[21]), .Z(n895) );
  OAI22_X2 U365 ( .A1(n898), .A2(n899), .B1(n394), .B2(n900), .ZN(n864) );
  NAND2_X2 U366 ( .A1(n869), .A2(n393), .ZN(n897) );
  NOR2_X2 U367 ( .A1(n1110), .A2(n901), .ZN(U7_Z_13) );
  XOR2_X2 U368 ( .A(n902), .B(n903), .Z(n901) );
  NAND2_X2 U371 ( .A1(n898), .A2(n899), .ZN(n869) );
  XOR2_X2 U372 ( .A(n905), .B(n906), .Z(n899) );
  NOR2_X2 U375 ( .A1(n893), .A2(in4[13]), .ZN(n841) );
  XOR2_X2 U376 ( .A(in2[31]), .B(n907), .Z(n893) );
  XOR2_X2 U377 ( .A(in2[20]), .B(in2[16]), .Z(n907) );
  XNOR2_X2 U378 ( .A(n908), .B(n909), .ZN(n898) );
  NAND2_X2 U381 ( .A1(n888), .A2(n501), .ZN(n855) );
  XOR2_X2 U382 ( .A(n426), .B(in1[30]), .Z(n888) );
  NOR2_X2 U383 ( .A1(n1110), .A2(n911), .ZN(U7_Z_12) );
  XNOR2_X2 U384 ( .A(n896), .B(n912), .ZN(n911) );
  NAND2_X2 U385 ( .A1(n900), .A2(n393), .ZN(n912) );
  NOR2_X2 U386 ( .A1(n913), .A2(n914), .ZN(n904) );
  NAND2_X2 U387 ( .A1(n914), .A2(n913), .ZN(n900) );
  XOR2_X2 U388 ( .A(n886), .B(n915), .Z(n913) );
  NOR2_X2 U389 ( .A1(n910), .A2(n887), .ZN(n915) );
  NOR2_X2 U390 ( .A1(n916), .A2(in3[12]), .ZN(n910) );
  XOR2_X2 U391 ( .A(in1[29]), .B(n917), .Z(n916) );
  XOR2_X2 U392 ( .A(in1[22]), .B(in1[31]), .Z(n917) );
  NAND2_X2 U393 ( .A1(n401), .A2(n918), .ZN(n886) );
  NAND3_X2 U394 ( .A1(n854), .A2(n402), .A3(n853), .ZN(n918) );
  OAI221_X2 U395 ( .B1(n919), .B2(n920), .C1(n409), .C2(n921), .A(n922), .ZN(
        n849) );
  NAND2_X2 U396 ( .A1(n923), .A2(n402), .ZN(n921) );
  XOR2_X2 U397 ( .A(n892), .B(n925), .Z(n914) );
  NOR2_X2 U398 ( .A1(n842), .A2(n894), .ZN(n925) );
  NOR2_X2 U399 ( .A1(n926), .A2(in4[12]), .ZN(n842) );
  XNOR2_X2 U400 ( .A(n463), .B(n927), .ZN(n926) );
  XOR2_X2 U401 ( .A(in2[19]), .B(in2[15]), .Z(n927) );
  NAND2_X2 U402 ( .A1(n832), .A2(n928), .ZN(n892) );
  NAND3_X2 U403 ( .A1(n839), .A2(n840), .A3(n838), .ZN(n928) );
  NOR2_X2 U406 ( .A1(n1110), .A2(n939), .ZN(U7_Z_11) );
  XOR2_X2 U407 ( .A(n940), .B(n941), .Z(n939) );
  NAND2_X2 U409 ( .A1(n942), .A2(n943), .ZN(n936) );
  NOR2_X2 U410 ( .A1(n943), .A2(n942), .ZN(n867) );
  XOR2_X2 U411 ( .A(n944), .B(n945), .Z(n942) );
  AOI221_X2 U412 ( .B1(n838), .B2(n839), .C1(n929), .C2(n932), .A(n471), .ZN(
        n945) );
  AND3_X2 U413 ( .A1(n932), .A2(n477), .A3(n947), .ZN(n838) );
  NAND2_X2 U414 ( .A1(n840), .A2(n931), .ZN(n944) );
  NAND2_X2 U415 ( .A1(in4[11]), .A2(n948), .ZN(n931) );
  XOR2_X2 U416 ( .A(in2[29]), .B(n949), .Z(n948) );
  XOR2_X2 U417 ( .A(in2[18]), .B(in2[14]), .Z(n949) );
  XOR2_X2 U418 ( .A(n950), .B(n951), .Z(n943) );
  AND3_X2 U420 ( .A1(n923), .A2(n413), .A3(n952), .ZN(n853) );
  NAND2_X2 U421 ( .A1(n402), .A2(n922), .ZN(n950) );
  NAND2_X2 U422 ( .A1(in3[11]), .A2(n953), .ZN(n922) );
  NOR2_X2 U423 ( .A1(n953), .A2(in3[11]), .ZN(n919) );
  XOR2_X2 U424 ( .A(in1[28]), .B(n954), .Z(n953) );
  XOR2_X2 U425 ( .A(in1[21]), .B(in1[30]), .Z(n954) );
  OAI221_X2 U426 ( .B1(n404), .B2(n938), .C1(n417), .C2(n866), .A(n935), .ZN(
        n940) );
  NAND3_X2 U427 ( .A1(n955), .A2(n510), .A3(n408), .ZN(n866) );
  NOR2_X2 U428 ( .A1(n1110), .A2(n956), .ZN(U7_Z_10) );
  XOR2_X2 U429 ( .A(n957), .B(n958), .Z(n956) );
  NAND2_X2 U430 ( .A1(n935), .A2(n955), .ZN(n958) );
  NAND2_X2 U431 ( .A1(n959), .A2(n960), .ZN(n955) );
  XNOR2_X2 U432 ( .A(n961), .B(n962), .ZN(n959) );
  OAI22_X2 U434 ( .A1(n964), .A2(n502), .B1(n410), .B2(n965), .ZN(n924) );
  NOR2_X2 U435 ( .A1(n966), .A2(n410), .ZN(n963) );
  NAND2_X2 U436 ( .A1(n920), .A2(n923), .ZN(n961) );
  NAND2_X2 U437 ( .A1(in3[10]), .A2(n967), .ZN(n920) );
  XOR2_X2 U438 ( .A(in1[27]), .B(n968), .Z(n967) );
  XOR2_X2 U439 ( .A(in1[20]), .B(in1[29]), .Z(n968) );
  XNOR2_X2 U440 ( .A(n969), .B(n970), .ZN(n960) );
  OAI22_X2 U442 ( .A1(n972), .A2(n505), .B1(n474), .B2(n973), .ZN(n929) );
  NOR2_X2 U443 ( .A1(n974), .A2(n474), .ZN(n971) );
  NAND2_X2 U444 ( .A1(n946), .A2(n932), .ZN(n969) );
  NAND2_X2 U445 ( .A1(in4[10]), .A2(n975), .ZN(n946) );
  XOR2_X2 U446 ( .A(in2[28]), .B(n976), .Z(n975) );
  XOR2_X2 U447 ( .A(in2[17]), .B(in2[13]), .Z(n976) );
  NOR2_X2 U450 ( .A1(n978), .A2(n979), .ZN(n511) );
  NAND2_X2 U451 ( .A1(n408), .A2(n510), .ZN(n977) );
  NAND2_X2 U452 ( .A1(n979), .A2(n978), .ZN(n510) );
  XNOR2_X2 U453 ( .A(n854), .B(n980), .ZN(n978) );
  NOR2_X2 U454 ( .A1(n415), .A2(n966), .ZN(n980) );
  XNOR2_X2 U455 ( .A(n839), .B(n981), .ZN(n979) );
  NOR2_X2 U456 ( .A1(n478), .A2(n974), .ZN(n981) );
  NOR2_X2 U457 ( .A1(n513), .A2(n512), .ZN(n514) );
  XOR2_X2 U458 ( .A(n982), .B(n983), .Z(n512) );
  NAND2_X2 U460 ( .A1(in3[8]), .A2(n984), .ZN(n965) );
  NOR2_X2 U461 ( .A1(n984), .A2(in3[8]), .ZN(n966) );
  XNOR2_X2 U462 ( .A(n420), .B(n985), .ZN(n984) );
  XOR2_X2 U463 ( .A(in1[18]), .B(in1[27]), .Z(n985) );
  NAND2_X2 U464 ( .A1(n986), .A2(n987), .ZN(n854) );
  NAND3_X2 U467 ( .A1(n424), .A2(n994), .A3(n421), .ZN(n992) );
  NAND2_X2 U469 ( .A1(n964), .A2(n502), .ZN(n952) );
  XNOR2_X2 U470 ( .A(in1[26]), .B(n995), .ZN(n964) );
  XOR2_X2 U471 ( .A(in1[19]), .B(in1[28]), .Z(n995) );
  XOR2_X2 U472 ( .A(n996), .B(n997), .Z(n513) );
  NAND2_X2 U474 ( .A1(in4[8]), .A2(n998), .ZN(n973) );
  NOR2_X2 U475 ( .A1(n998), .A2(in4[8]), .ZN(n974) );
  XOR2_X2 U476 ( .A(in2[11]), .B(n999), .Z(n998) );
  XOR2_X2 U477 ( .A(in2[26]), .B(in2[15]), .Z(n999) );
  NAND2_X2 U478 ( .A1(n1000), .A2(n1001), .ZN(n839) );
  NAND3_X2 U481 ( .A1(n488), .A2(n1008), .A3(n486), .ZN(n1006) );
  NAND2_X2 U483 ( .A1(n972), .A2(n505), .ZN(n947) );
  XNOR2_X2 U484 ( .A(in2[12]), .B(n1009), .ZN(n972) );
  XOR2_X2 U485 ( .A(in2[27]), .B(in2[16]), .Z(n1009) );
  NAND2_X2 U486 ( .A1(n521), .A2(n1010), .ZN(n509) );
  NAND2_X2 U488 ( .A1(n1012), .A2(n1013), .ZN(n520) );
  NOR2_X2 U489 ( .A1(n1014), .A2(n1015), .ZN(n524) );
  NAND2_X2 U491 ( .A1(n1015), .A2(n1014), .ZN(n523) );
  XNOR2_X2 U492 ( .A(n1017), .B(n1018), .ZN(n1014) );
  NOR2_X2 U493 ( .A1(n1003), .A2(n1007), .ZN(n1018) );
  XNOR2_X2 U494 ( .A(n1019), .B(n1020), .ZN(n1015) );
  NOR2_X2 U495 ( .A1(n989), .A2(n993), .ZN(n1020) );
  NAND3_X2 U496 ( .A1(n533), .A2(n532), .A3(n536), .ZN(n1016) );
  NAND2_X2 U501 ( .A1(n1027), .A2(n1028), .ZN(n588) );
  NAND2_X2 U502 ( .A1(n592), .A2(n593), .ZN(n591) );
  XOR2_X2 U503 ( .A(n492), .B(n1029), .Z(n593) );
  XOR2_X2 U505 ( .A(n1032), .B(n1033), .Z(n592) );
  NOR2_X2 U507 ( .A1(n1028), .A2(n1027), .ZN(n1021) );
  XOR2_X2 U508 ( .A(n1036), .B(n1037), .Z(n1027) );
  NOR2_X2 U510 ( .A1(in4[2]), .A2(n1030), .ZN(n1039) );
  XOR2_X2 U511 ( .A(n1041), .B(n1042), .Z(n1028) );
  NOR2_X2 U513 ( .A1(in3[2]), .A2(n1034), .ZN(n1044) );
  NAND2_X2 U514 ( .A1(n1045), .A2(n1046), .ZN(n533) );
  OAI22_X2 U515 ( .A1(n534), .A2(n535), .B1(n423), .B2(n531), .ZN(n1047) );
  XNOR2_X2 U516 ( .A(n994), .B(n1048), .ZN(n1045) );
  NOR2_X2 U517 ( .A1(n1049), .A2(n425), .ZN(n1048) );
  XNOR2_X2 U518 ( .A(n1008), .B(n1050), .ZN(n1046) );
  NOR2_X2 U519 ( .A1(n1051), .A2(n489), .ZN(n1050) );
  NAND2_X2 U520 ( .A1(n534), .A2(n535), .ZN(n536) );
  XNOR2_X2 U521 ( .A(n1052), .B(n1053), .ZN(n535) );
  NAND2_X2 U523 ( .A1(n1056), .A2(n1057), .ZN(n1052) );
  XNOR2_X2 U524 ( .A(n1058), .B(n1059), .ZN(n534) );
  NAND2_X2 U526 ( .A1(n1062), .A2(n1063), .ZN(n1058) );
  XNOR2_X2 U527 ( .A(n1064), .B(n1065), .ZN(n1012) );
  NAND2_X2 U531 ( .A1(in4[4]), .A2(n1067), .ZN(n1062) );
  NAND2_X2 U532 ( .A1(n1008), .A2(n488), .ZN(n1063) );
  NOR2_X2 U533 ( .A1(n1067), .A2(in4[4]), .ZN(n1051) );
  XOR2_X2 U534 ( .A(in2[11]), .B(n1068), .Z(n1067) );
  XOR2_X2 U535 ( .A(in2[7]), .B(in2[22]), .Z(n1068) );
  NAND2_X2 U540 ( .A1(in4[3]), .A2(n1074), .ZN(n1038) );
  NAND2_X2 U541 ( .A1(in4[2]), .A2(n1030), .ZN(n1031) );
  XOR2_X2 U542 ( .A(in2[20]), .B(n1075), .Z(n1030) );
  XOR2_X2 U543 ( .A(in2[9]), .B(in2[5]), .Z(n1075) );
  NOR2_X2 U544 ( .A1(n1074), .A2(in4[3]), .ZN(n1069) );
  XOR2_X2 U545 ( .A(in2[10]), .B(n1076), .Z(n1074) );
  XOR2_X2 U546 ( .A(in2[6]), .B(in2[21]), .Z(n1076) );
  NOR2_X2 U547 ( .A1(n1060), .A2(in4[5]), .ZN(n1061) );
  XOR2_X2 U548 ( .A(in2[12]), .B(n1077), .Z(n1060) );
  XOR2_X2 U549 ( .A(in2[8]), .B(in2[23]), .Z(n1077) );
  NOR2_X2 U550 ( .A1(n1066), .A2(in4[6]), .ZN(n1007) );
  XOR2_X2 U551 ( .A(in2[13]), .B(n1078), .Z(n1066) );
  XOR2_X2 U552 ( .A(in2[9]), .B(in2[24]), .Z(n1078) );
  NAND2_X2 U553 ( .A1(n1004), .A2(n1000), .ZN(n1064) );
  NAND2_X2 U554 ( .A1(in4[7]), .A2(n1079), .ZN(n1000) );
  XOR2_X2 U555 ( .A(in2[10]), .B(n1080), .Z(n1079) );
  XOR2_X2 U556 ( .A(in2[25]), .B(in2[14]), .Z(n1080) );
  XNOR2_X2 U557 ( .A(n1081), .B(n1082), .ZN(n1013) );
  NAND2_X2 U561 ( .A1(in3[4]), .A2(n1084), .ZN(n1056) );
  NAND2_X2 U562 ( .A1(n994), .A2(n424), .ZN(n1057) );
  NOR2_X2 U563 ( .A1(n1084), .A2(in3[4]), .ZN(n1049) );
  XNOR2_X2 U564 ( .A(n1085), .B(in1[14]), .ZN(n1084) );
  XOR2_X2 U565 ( .A(in1[21]), .B(n426), .Z(n1085) );
  NAND2_X2 U569 ( .A1(n1089), .A2(n1090), .ZN(n1088) );
  NAND2_X2 U570 ( .A1(in3[3]), .A2(n1091), .ZN(n1043) );
  NAND2_X2 U571 ( .A1(in3[2]), .A2(n1034), .ZN(n1035) );
  XNOR2_X2 U572 ( .A(n1092), .B(in1[12]), .ZN(n1034) );
  XNOR2_X2 U573 ( .A(in1[19]), .B(in1[21]), .ZN(n1092) );
  NOR2_X2 U574 ( .A1(n1091), .A2(in3[3]), .ZN(n1086) );
  XNOR2_X2 U575 ( .A(n1093), .B(in1[13]), .ZN(n1091) );
  XNOR2_X2 U576 ( .A(in1[20]), .B(in1[22]), .ZN(n1093) );
  NOR2_X2 U577 ( .A1(n1054), .A2(in3[5]), .ZN(n1055) );
  XNOR2_X2 U578 ( .A(n1094), .B(in1[15]), .ZN(n1054) );
  XNOR2_X2 U579 ( .A(in1[22]), .B(in1[24]), .ZN(n1094) );
  NOR2_X2 U580 ( .A1(n1083), .A2(in3[6]), .ZN(n993) );
  XNOR2_X2 U581 ( .A(n420), .B(n1095), .ZN(n1083) );
  XOR2_X2 U582 ( .A(in1[23]), .B(in1[16]), .Z(n1095) );
  NAND2_X2 U583 ( .A1(n990), .A2(n986), .ZN(n1081) );
  NAND2_X2 U584 ( .A1(in3[7]), .A2(n1096), .ZN(n986) );
  XOR2_X2 U585 ( .A(in1[26]), .B(n1097), .Z(n1096) );
  XOR2_X2 U586 ( .A(in1[24]), .B(in1[17]), .Z(n1097) );
  NOR2_X2 U587 ( .A1(n1110), .A2(n1098), .ZN(U7_Z_1) );
  XNOR2_X2 U588 ( .A(n1026), .B(n1099), .ZN(n1098) );
  XOR2_X2 U589 ( .A(n1024), .B(n1023), .Z(n1099) );
  XNOR2_X2 U590 ( .A(n1071), .B(n1100), .ZN(n1023) );
  XOR2_X2 U591 ( .A(in4[1]), .B(n495), .Z(n1100) );
  XNOR2_X2 U592 ( .A(in2[19]), .B(n1101), .ZN(n1071) );
  XOR2_X2 U593 ( .A(in2[8]), .B(in2[4]), .Z(n1101) );
  XNOR2_X2 U594 ( .A(n1090), .B(n1102), .ZN(n1026) );
  XOR2_X2 U595 ( .A(in3[1]), .B(n433), .Z(n1102) );
  XOR2_X2 U596 ( .A(n1103), .B(in1[11]), .Z(n1090) );
  XNOR2_X2 U597 ( .A(in1[18]), .B(in1[20]), .ZN(n1103) );
  NOR2_X2 U599 ( .A1(n1105), .A2(n1104), .ZN(n1024) );
  NAND2_X2 U601 ( .A1(in3[0]), .A2(n1106), .ZN(n1089) );
  XNOR2_X2 U602 ( .A(n1107), .B(in1[10]), .ZN(n1106) );
  XNOR2_X2 U603 ( .A(in1[17]), .B(in1[19]), .ZN(n1107) );
  NAND2_X2 U605 ( .A1(in4[0]), .A2(n1108), .ZN(n1072) );
  XOR2_X2 U606 ( .A(in2[18]), .B(n1109), .Z(n1108) );
  XOR2_X2 U607 ( .A(in2[7]), .B(in2[3]), .Z(n1109) );
  INV_X4 U608 ( .A(n699), .ZN(n366) );
  INV_X4 U610 ( .A(n691), .ZN(n368) );
  INV_X4 U612 ( .A(n627), .ZN(n370) );
  INV_X4 U613 ( .A(n631), .ZN(n371) );
  INV_X4 U615 ( .A(n562), .ZN(n373) );
  INV_X4 U616 ( .A(n580), .ZN(n374) );
  INV_X4 U617 ( .A(n665), .ZN(n375) );
  INV_X4 U618 ( .A(n657), .ZN(n376) );
  INV_X4 U619 ( .A(n689), .ZN(n377) );
  INV_X4 U620 ( .A(n700), .ZN(n378) );
  INV_X4 U621 ( .A(n696), .ZN(n379) );
  INV_X4 U622 ( .A(n721), .ZN(n380) );
  INV_X4 U623 ( .A(n764), .ZN(n381) );
  INV_X4 U624 ( .A(n862), .ZN(n382) );
  INV_X4 U627 ( .A(n813), .ZN(n385) );
  INV_X4 U628 ( .A(n791), .ZN(n386) );
  INV_X4 U629 ( .A(n767), .ZN(n387) );
  INV_X4 U630 ( .A(n694), .ZN(n388) );
  INV_X4 U631 ( .A(n734), .ZN(n389) );
  INV_X4 U632 ( .A(n850), .ZN(n390) );
  INV_X4 U634 ( .A(n864), .ZN(n392) );
  INV_X4 U635 ( .A(n904), .ZN(n393) );
  INV_X4 U636 ( .A(n869), .ZN(n394) );
  INV_X4 U637 ( .A(n910), .ZN(n395) );
  INV_X4 U638 ( .A(n740), .ZN(n396) );
  INV_X4 U639 ( .A(n720), .ZN(n397) );
  INV_X4 U640 ( .A(n888), .ZN(n398) );
  INV_X4 U642 ( .A(n934), .ZN(n400) );
  INV_X4 U643 ( .A(n849), .ZN(n401) );
  INV_X4 U644 ( .A(n919), .ZN(n402) );
  INV_X4 U645 ( .A(n758), .ZN(n403) );
  INV_X4 U646 ( .A(n955), .ZN(n404) );
  INV_X4 U648 ( .A(n759), .ZN(n406) );
  INV_X4 U649 ( .A(n782), .ZN(n407) );
  INV_X4 U650 ( .A(n514), .ZN(n408) );
  INV_X4 U651 ( .A(n924), .ZN(n409) );
  INV_X4 U652 ( .A(n952), .ZN(n410) );
  INV_X4 U653 ( .A(n760), .ZN(n411) );
  INV_X4 U654 ( .A(n784), .ZN(n412) );
  INV_X4 U655 ( .A(n966), .ZN(n413) );
  INV_X4 U657 ( .A(n965), .ZN(n415) );
  INV_X4 U658 ( .A(n783), .ZN(n416) );
  INV_X4 U659 ( .A(n509), .ZN(n417) );
  INV_X4 U660 ( .A(n993), .ZN(n418) );
  INV_X4 U661 ( .A(n523), .ZN(n419) );
  INV_X4 U662 ( .A(in1[25]), .ZN(n420) );
  INV_X4 U663 ( .A(n1055), .ZN(n421) );
  INV_X4 U664 ( .A(n1047), .ZN(n422) );
  INV_X4 U665 ( .A(n536), .ZN(n423) );
  INV_X4 U666 ( .A(n1049), .ZN(n424) );
  INV_X4 U667 ( .A(n1056), .ZN(n425) );
  INV_X4 U668 ( .A(in1[23]), .ZN(n426) );
  INV_X4 U669 ( .A(n1021), .ZN(n427) );
  INV_X4 U670 ( .A(n1086), .ZN(n428) );
  INV_X4 U671 ( .A(n589), .ZN(n429) );
  INV_X4 U672 ( .A(n1025), .ZN(n430) );
  INV_X4 U673 ( .A(n1032), .ZN(n431) );
  INV_X4 U674 ( .A(n1090), .ZN(n432) );
  INV_X4 U675 ( .A(n1089), .ZN(n433) );
  INV_X4 U676 ( .A(in1[8]), .ZN(n434) );
  INV_X4 U677 ( .A(n554), .ZN(n435) );
  INV_X4 U678 ( .A(in1[7]), .ZN(n436) );
  INV_X4 U679 ( .A(n599), .ZN(n437) );
  INV_X4 U680 ( .A(in1[5]), .ZN(n438) );
  INV_X4 U681 ( .A(n643), .ZN(n439) );
  INV_X4 U682 ( .A(n615), .ZN(n440) );
  INV_X4 U683 ( .A(n619), .ZN(n441) );
  INV_X4 U684 ( .A(n621), .ZN(n442) );
  INV_X4 U685 ( .A(n620), .ZN(n443) );
  INV_X4 U686 ( .A(n666), .ZN(n444) );
  INV_X4 U687 ( .A(in1[1]), .ZN(n445) );
  INV_X4 U688 ( .A(n713), .ZN(n446) );
  INV_X4 U689 ( .A(n548), .ZN(n447) );
  INV_X4 U690 ( .A(n551), .ZN(n448) );
  INV_X4 U691 ( .A(n552), .ZN(n449) );
  INV_X4 U692 ( .A(n624), .ZN(n450) );
  INV_X4 U693 ( .A(n611), .ZN(n451) );
  INV_X4 U694 ( .A(n652), .ZN(n452) );
  INV_X4 U695 ( .A(n612), .ZN(n453) );
  INV_X4 U696 ( .A(n861), .ZN(n454) );
  INV_X4 U697 ( .A(n692), .ZN(n455) );
  INV_X4 U698 ( .A(n672), .ZN(n456) );
  INV_X4 U699 ( .A(n827), .ZN(n457) );
  INV_X4 U700 ( .A(n834), .ZN(n458) );
  INV_X4 U701 ( .A(n841), .ZN(n459) );
  INV_X4 U702 ( .A(n833), .ZN(n460) );
  INV_X4 U703 ( .A(n680), .ZN(n461) );
  INV_X4 U704 ( .A(n842), .ZN(n462) );
  INV_X4 U705 ( .A(in2[30]), .ZN(n463) );
  INV_X4 U706 ( .A(n638), .ZN(n464) );
  INV_X4 U707 ( .A(n607), .ZN(n465) );
  INV_X4 U708 ( .A(n709), .ZN(n466) );
  INV_X4 U710 ( .A(n613), .ZN(n468) );
  INV_X4 U711 ( .A(n679), .ZN(n469) );
  INV_X4 U712 ( .A(n727), .ZN(n470) );
  INV_X4 U713 ( .A(n946), .ZN(n471) );
  INV_X4 U714 ( .A(n726), .ZN(n472) );
  INV_X4 U715 ( .A(n737), .ZN(n473) );
  INV_X4 U716 ( .A(n947), .ZN(n474) );
  INV_X4 U717 ( .A(n748), .ZN(n475) );
  INV_X4 U718 ( .A(in2[26]), .ZN(n476) );
  INV_X4 U719 ( .A(n974), .ZN(n477) );
  INV_X4 U720 ( .A(n973), .ZN(n478) );
  INV_X4 U721 ( .A(n788), .ZN(n479) );
  INV_X4 U722 ( .A(n749), .ZN(n480) );
  INV_X4 U723 ( .A(n787), .ZN(n481) );
  INV_X4 U724 ( .A(n802), .ZN(n482) );
  INV_X4 U725 ( .A(n1007), .ZN(n483) );
  INV_X4 U726 ( .A(n804), .ZN(n484) );
  INV_X4 U727 ( .A(n789), .ZN(n485) );
  INV_X4 U728 ( .A(n1061), .ZN(n486) );
  INV_X4 U730 ( .A(n1051), .ZN(n488) );
  INV_X4 U731 ( .A(n1062), .ZN(n489) );
  INV_X4 U733 ( .A(n1069), .ZN(n491) );
  INV_X4 U734 ( .A(n1040), .ZN(n492) );
  INV_X4 U735 ( .A(n1071), .ZN(n493) );
  INV_X4 U737 ( .A(n1072), .ZN(n495) );
  INV_X4 U738 ( .A(n549), .ZN(n496) );
  INV_X4 U739 ( .A(in3[30]), .ZN(n497) );
  INV_X4 U740 ( .A(in3[29]), .ZN(n498) );
  INV_X4 U741 ( .A(in3[23]), .ZN(n499) );
  INV_X4 U742 ( .A(in3[15]), .ZN(n500) );
  INV_X4 U743 ( .A(in3[13]), .ZN(n501) );
  INV_X4 U744 ( .A(in3[9]), .ZN(n502) );
  INV_X4 U745 ( .A(in4[23]), .ZN(n503) );
  INV_X4 U746 ( .A(in4[17]), .ZN(n504) );
  INV_X4 U747 ( .A(in4[9]), .ZN(n505) );
  OR2_X1 U748 ( .A1(n419), .A2(n524), .ZN(n526) );
  AND2_X1 U749 ( .A1(n437), .A2(n558), .ZN(n583) );
  AND2_X1 U750 ( .A1(in4[28]), .A2(in2[31]), .ZN(n575) );
  AND2_X1 U751 ( .A1(in3[28]), .A2(in1[6]), .ZN(n584) );
  OR2_X1 U752 ( .A1(n376), .A2(n630), .ZN(n653) );
  OR2_X1 U753 ( .A1(in1[0]), .A2(in3[22]), .ZN(n686) );
  AND2_X1 U754 ( .A1(in4[22]), .A2(n723), .ZN(n678) );
  AND2_X1 U755 ( .A1(n752), .A2(n475), .ZN(n746) );
  AND2_X1 U756 ( .A1(n763), .A2(n403), .ZN(n756) );
  AND2_X1 U757 ( .A1(in3[16]), .A2(in1[26]), .ZN(n808) );
  OR4_X1 U758 ( .A1(n866), .A2(n856), .A3(n417), .A4(n867), .ZN(n857) );
  AND2_X1 U759 ( .A1(n851), .A2(n885), .ZN(n879) );
  AND2_X1 U760 ( .A1(n836), .A2(n891), .ZN(n876) );
  AND2_X1 U761 ( .A1(in3[12]), .A2(n916), .ZN(n887) );
  AND2_X1 U762 ( .A1(in4[12]), .A2(n926), .ZN(n894) );
  AND2_X1 U763 ( .A1(n932), .A2(n840), .ZN(n930) );
  AND2_X1 U764 ( .A1(n400), .A2(n933), .ZN(n896) );
  OR3_X1 U765 ( .A1(n417), .A2(n867), .A3(n866), .ZN(n933) );
  OR3_X1 U766 ( .A1(n404), .A2(n867), .A3(n938), .ZN(n937) );
  OR2_X1 U767 ( .A1(n948), .A2(in4[11]), .ZN(n840) );
  OR2_X1 U768 ( .A1(n960), .A2(n959), .ZN(n935) );
  OR2_X1 U769 ( .A1(n967), .A2(in3[10]), .ZN(n923) );
  OR2_X1 U770 ( .A1(n975), .A2(in4[10]), .ZN(n932) );
  AND2_X1 U771 ( .A1(n1038), .A2(n491), .ZN(n1037) );
  AND2_X1 U772 ( .A1(n1043), .A2(n428), .ZN(n1042) );
  OR2_X1 U773 ( .A1(n1046), .A2(n1045), .ZN(n531) );
  OR2_X1 U774 ( .A1(n1013), .A2(n1012), .ZN(n521) );
  AND2_X1 U775 ( .A1(in4[6]), .A2(n1066), .ZN(n1003) );
  OR2_X1 U776 ( .A1(n1079), .A2(in4[7]), .ZN(n1004) );
  AND2_X1 U777 ( .A1(in3[6]), .A2(n1083), .ZN(n989) );
  OR2_X1 U778 ( .A1(n1096), .A2(in3[7]), .ZN(n990) );
  DFF_X2 ops_out_reg_0_ ( .D(U7_Z_0), .CK(clock), .Q(ops_out[0]) );
  DFF_X2 ops_out_reg_1_ ( .D(U7_Z_1), .CK(clock), .Q(ops_out[1]) );
  DFF_X2 ops_out_reg_2_ ( .D(U7_Z_2), .CK(clock), .Q(ops_out[2]) );
  DFF_X2 ops_out_reg_3_ ( .D(U7_Z_3), .CK(clock), .Q(ops_out[3]) );
  DFF_X2 ops_out_reg_4_ ( .D(U7_Z_4), .CK(clock), .Q(ops_out[4]) );
  DFF_X2 ops_out_reg_5_ ( .D(U7_Z_5), .CK(clock), .Q(ops_out[5]) );
  DFF_X2 ops_out_reg_6_ ( .D(U7_Z_6), .CK(clock), .Q(ops_out[6]) );
  DFF_X2 ops_out_reg_7_ ( .D(U7_Z_7), .CK(clock), .Q(ops_out[7]) );
  DFF_X2 ops_out_reg_8_ ( .D(U7_Z_8), .CK(clock), .Q(ops_out[8]) );
  DFF_X2 ops_out_reg_9_ ( .D(U7_Z_9), .CK(clock), .Q(ops_out[9]) );
  DFF_X2 ops_out_reg_10_ ( .D(U7_Z_10), .CK(clock), .Q(ops_out[10]) );
  DFF_X2 ops_out_reg_11_ ( .D(U7_Z_11), .CK(clock), .Q(ops_out[11]) );
  DFF_X2 ops_out_reg_12_ ( .D(U7_Z_12), .CK(clock), .Q(ops_out[12]) );
  DFF_X2 ops_out_reg_13_ ( .D(U7_Z_13), .CK(clock), .Q(ops_out[13]) );
  DFF_X2 ops_out_reg_14_ ( .D(U7_Z_14), .CK(clock), .Q(ops_out[14]) );
  DFF_X2 ops_out_reg_15_ ( .D(U7_Z_15), .CK(clock), .Q(ops_out[15]) );
  DFF_X2 ops_out_reg_16_ ( .D(U7_Z_16), .CK(clock), .Q(ops_out[16]) );
  DFF_X2 ops_out_reg_17_ ( .D(U7_Z_17), .CK(clock), .Q(ops_out[17]) );
  DFF_X2 ops_out_reg_18_ ( .D(U7_Z_18), .CK(clock), .Q(ops_out[18]) );
  DFF_X2 ops_out_reg_19_ ( .D(U7_Z_19), .CK(clock), .Q(ops_out[19]) );
  DFF_X2 ops_out_reg_20_ ( .D(U7_Z_20), .CK(clock), .Q(ops_out[20]) );
  DFF_X2 ops_out_reg_21_ ( .D(U7_Z_21), .CK(clock), .Q(ops_out[21]) );
  DFF_X2 ops_out_reg_22_ ( .D(U7_Z_22), .CK(clock), .Q(ops_out[22]) );
  DFF_X2 ops_out_reg_23_ ( .D(U7_Z_23), .CK(clock), .Q(ops_out[23]) );
  DFF_X2 ops_out_reg_24_ ( .D(U7_Z_24), .CK(clock), .Q(ops_out[24]) );
  DFF_X2 ops_out_reg_25_ ( .D(U7_Z_25), .CK(clock), .Q(ops_out[25]) );
  DFF_X2 ops_out_reg_26_ ( .D(U7_Z_26), .CK(clock), .Q(ops_out[26]) );
  DFF_X2 ops_out_reg_27_ ( .D(U7_Z_27), .CK(clock), .Q(ops_out[27]) );
  DFF_X2 ops_out_reg_28_ ( .D(U7_Z_28), .CK(clock), .Q(ops_out[28]) );
  DFF_X2 ops_out_reg_29_ ( .D(U7_Z_29), .CK(clock), .Q(ops_out[29]) );
  DFF_X2 ops_out_reg_30_ ( .D(U7_Z_30), .CK(clock), .Q(ops_out[30]) );
  DFF_X2 ops_out_reg_31_ ( .D(U7_Z_31), .CK(clock), .Q(ops_out[31]) );
  OR2_X4 U779 ( .A1(n861), .A2(n859), .ZN(n868) );
  AOI222_X1 U780 ( .A1(n929), .A2(n930), .B1(in4[11]), .B2(n948), .C1(n471), 
        .C2(n840), .ZN(n832) );
  AOI222_X1 U781 ( .A1(in3[10]), .A2(n967), .B1(n854), .B2(n853), .C1(n923), 
        .C2(n924), .ZN(n951) );
  XOR2_X2 U782 ( .A(in2[22]), .B(in2[26]), .Z(n790) );
  OAI21_X2 U783 ( .B1(n895), .B2(in4[14]), .A(n837), .ZN(n890) );
  OAI21_X2 U784 ( .B1(n943), .B2(n942), .A(n936), .ZN(n941) );
  XOR2_X2 U785 ( .A(in2[18]), .B(in2[22]), .Z(n828) );
  OAI21_X2 U786 ( .B1(n604), .B2(n605), .A(n566), .ZN(n603) );
  AOI21_X2 U787 ( .B1(n669), .B2(n670), .A(n630), .ZN(n668) );
  OAI21_X2 U788 ( .B1(n716), .B2(n717), .A(n695), .ZN(n715) );
  OAI21_X2 U789 ( .B1(n823), .B2(n824), .A(n792), .ZN(n822) );
  OAI21_X2 U790 ( .B1(n882), .B2(n883), .A(n863), .ZN(n881) );
  OAI21_X2 U791 ( .B1(n978), .B2(n979), .A(n510), .ZN(n516) );
  OAI211_X2 U792 ( .C1(n867), .C2(n935), .A(n936), .B(n937), .ZN(n934) );
  AOI21_X2 U793 ( .B1(n764), .B2(n765), .A(n766), .ZN(n698) );
  AOI22_X2 U794 ( .A1(n513), .A2(n512), .B1(n408), .B2(n511), .ZN(n938) );
  AOI21_X2 U795 ( .B1(n863), .B2(n864), .A(n865), .ZN(n862) );
  OAI21_X2 U796 ( .B1(n1011), .B2(n524), .A(n520), .ZN(n1010) );
  AOI21_X2 U797 ( .B1(n422), .B2(n1016), .A(n419), .ZN(n1011) );
  OAI21_X2 U798 ( .B1(n629), .B2(n653), .A(n370), .ZN(n639) );
  AOI21_X2 U799 ( .B1(n695), .B2(n700), .A(n701), .ZN(n699) );
  OAI21_X2 U800 ( .B1(n698), .B2(n728), .A(n378), .ZN(n705) );
  OAI21_X2 U801 ( .B1(n896), .B2(n897), .A(n392), .ZN(n873) );
  OAI21_X2 U802 ( .B1(n417), .B2(n977), .A(n938), .ZN(n957) );
  OAI21_X2 U803 ( .B1(n423), .B2(n527), .A(n422), .ZN(n522) );
  AOI21_X2 U804 ( .B1(n509), .B2(n510), .A(n511), .ZN(n508) );
  AOI21_X2 U805 ( .B1(n512), .B2(n513), .A(n514), .ZN(n507) );
  AOI21_X2 U806 ( .B1(n522), .B2(n523), .A(n524), .ZN(n518) );
  OAI21_X2 U807 ( .B1(n589), .B2(n590), .A(n591), .ZN(n586) );
  OAI211_X2 U808 ( .C1(n450), .C2(n371), .A(n622), .B(n623), .ZN(n564) );
  OAI21_X2 U809 ( .B1(n631), .B2(n624), .A(n625), .ZN(n622) );
  OAI21_X2 U810 ( .B1(n964), .B2(n502), .A(n952), .ZN(n982) );
  AOI21_X2 U811 ( .B1(n854), .B2(n413), .A(n415), .ZN(n983) );
  OAI21_X2 U812 ( .B1(n803), .B2(n504), .A(n802), .ZN(n819) );
  AOI21_X2 U813 ( .B1(n485), .B2(n457), .A(n484), .ZN(n820) );
  OAI21_X2 U814 ( .B1(n420), .B2(n500), .A(n847), .ZN(n877) );
  OAI21_X2 U815 ( .B1(n879), .B2(n850), .A(n852), .ZN(n878) );
  OAI21_X2 U816 ( .B1(n988), .B2(n989), .A(n990), .ZN(n987) );
  AOI21_X2 U817 ( .B1(n991), .B2(n992), .A(n993), .ZN(n988) );
  OAI211_X2 U818 ( .C1(n400), .C2(n856), .A(n857), .B(n858), .ZN(n764) );
  AOI22_X2 U819 ( .A1(n859), .A2(n860), .B1(n861), .B2(n382), .ZN(n858) );
  OAI211_X2 U820 ( .C1(n420), .C2(n500), .A(n844), .B(n845), .ZN(n755) );
  AOI22_X2 U821 ( .A1(n846), .A2(n847), .B1(n848), .B2(n849), .ZN(n845) );
  OAI21_X2 U822 ( .B1(n888), .B2(n501), .A(n855), .ZN(n908) );
  AOI21_X2 U823 ( .B1(n886), .B2(n395), .A(n887), .ZN(n909) );
  OAI21_X2 U824 ( .B1(n1002), .B2(n1003), .A(n1004), .ZN(n1001) );
  AOI21_X2 U825 ( .B1(n1005), .B2(n1006), .A(n1007), .ZN(n1002) );
  AOI22_X2 U826 ( .A1(n810), .A2(n811), .B1(n385), .B2(n812), .ZN(n769) );
  AOI21_X2 U827 ( .B1(n1023), .B2(n1024), .A(n430), .ZN(n589) );
  OAI21_X2 U828 ( .B1(n1024), .B2(n1023), .A(n1026), .ZN(n1025) );
  OAI211_X2 U829 ( .C1(n1021), .C2(n591), .A(n588), .B(n1022), .ZN(n532) );
  OAI211_X2 U830 ( .C1(n592), .C2(n593), .A(n429), .B(n427), .ZN(n1022) );
  OAI211_X2 U831 ( .C1(n559), .C2(n560), .A(n561), .B(n373), .ZN(n542) );
  AOI21_X2 U832 ( .B1(n560), .B2(n559), .A(n563), .ZN(n562) );
  OAI21_X2 U833 ( .B1(n972), .B2(n505), .A(n947), .ZN(n996) );
  AOI21_X2 U834 ( .B1(n839), .B2(n477), .A(n478), .ZN(n997) );
  AOI21_X2 U835 ( .B1(n368), .B2(n455), .A(n698), .ZN(n697) );
  AOI21_X2 U836 ( .B1(n628), .B2(n639), .A(n631), .ZN(n634) );
  AOI21_X2 U837 ( .B1(n578), .B2(n577), .A(n580), .ZN(n595) );
  AOI21_X2 U838 ( .B1(n564), .B2(n566), .A(n579), .ZN(n596) );
  OAI21_X2 U839 ( .B1(n436), .B2(n498), .A(n558), .ZN(n597) );
  AOI21_X2 U840 ( .B1(n556), .B2(n437), .A(n584), .ZN(n598) );
  OAI21_X2 U841 ( .B1(n674), .B2(n503), .A(n680), .ZN(n706) );
  AOI21_X2 U842 ( .B1(n708), .B2(n466), .A(n678), .ZN(n707) );
  AOI22_X2 U843 ( .A1(n577), .A2(n578), .B1(n374), .B2(n579), .ZN(n559) );
  AOI21_X2 U844 ( .B1(n457), .B2(n746), .A(n747), .ZN(n677) );
  AOI21_X2 U845 ( .B1(n755), .B2(n756), .A(n757), .ZN(n688) );
  OAI21_X2 U846 ( .B1(n688), .B2(n719), .A(n689), .ZN(n712) );
  AOI21_X2 U847 ( .B1(n705), .B2(n695), .A(n701), .ZN(n704) );
  OAI21_X2 U848 ( .B1(n677), .B2(n724), .A(n679), .ZN(n708) );
  OAI21_X2 U849 ( .B1(n456), .B2(n651), .A(n611), .ZN(n637) );
  OAI21_X2 U850 ( .B1(n375), .B2(n649), .A(n619), .ZN(n642) );
  OAI21_X2 U851 ( .B1(n1055), .B2(n1057), .A(n991), .ZN(n1019) );
  OAI21_X2 U852 ( .B1(n1061), .B2(n1063), .A(n1005), .ZN(n1017) );
  AOI21_X2 U853 ( .B1(n963), .B2(n854), .A(n924), .ZN(n962) );
  AOI21_X2 U854 ( .B1(n483), .B2(n1017), .A(n1003), .ZN(n1065) );
  AOI21_X2 U855 ( .B1(n971), .B2(n839), .A(n929), .ZN(n970) );
  AOI21_X2 U856 ( .B1(n418), .B2(n1019), .A(n989), .ZN(n1082) );
  OAI21_X2 U857 ( .B1(n850), .B2(n851), .A(n852), .ZN(n846) );
  OAI21_X2 U858 ( .B1(n835), .B2(n836), .A(n837), .ZN(n834) );
  OAI21_X2 U859 ( .B1(n654), .B2(n655), .A(n657), .ZN(n659) );
  OAI21_X2 U860 ( .B1(n630), .B2(n629), .A(n656), .ZN(n660) );
  AOI21_X2 U861 ( .B1(n469), .B2(n466), .A(n678), .ZN(n673) );
  AOI21_X2 U862 ( .B1(n811), .B2(n810), .A(n813), .ZN(n815) );
  AOI21_X2 U863 ( .B1(n792), .B2(n764), .A(n812), .ZN(n816) );
  OAI21_X2 U864 ( .B1(n898), .B2(n899), .A(n869), .ZN(n902) );
  OAI21_X2 U865 ( .B1(n904), .B2(n896), .A(n900), .ZN(n903) );
  OAI21_X2 U866 ( .B1(n729), .B2(n730), .A(n696), .ZN(n732) );
  OAI21_X2 U867 ( .B1(n388), .B2(n698), .A(n389), .ZN(n733) );
  AOI21_X2 U868 ( .B1(n873), .B2(n863), .A(n865), .ZN(n872) );
  OAI21_X2 U869 ( .B1(n534), .B2(n535), .A(n536), .ZN(n529) );
  OAI21_X2 U870 ( .B1(n592), .B2(n593), .A(n591), .ZN(n774) );
  AOI211_X2 U871 ( .C1(n1104), .C2(n1105), .A(n1110), .B(n1024), .ZN(U7_Z_0)
         );
  INV_X4 U872 ( .A(n1111), .ZN(n1110) );
  AOI21_X2 U873 ( .B1(in4[15]), .B2(n828), .A(n831), .ZN(n875) );
  OAI21_X2 U874 ( .B1(n835), .B2(n876), .A(n837), .ZN(n874) );
  AOI21_X2 U875 ( .B1(in1[27]), .B2(in3[17]), .A(n784), .ZN(n817) );
  AOI21_X2 U876 ( .B1(n416), .B2(n755), .A(n808), .ZN(n818) );
  AOI21_X2 U877 ( .B1(n893), .B2(in4[13]), .A(n841), .ZN(n905) );
  AOI21_X2 U878 ( .B1(n892), .B2(n462), .A(n894), .ZN(n906) );
  AOI22_X2 U879 ( .A1(n432), .A2(n433), .B1(n1088), .B2(in3[1]), .ZN(n1032) );
  AOI22_X2 U880 ( .A1(n1060), .A2(in4[5]), .B1(n486), .B2(n489), .ZN(n1005) );
  AOI21_X2 U881 ( .B1(in3[5]), .B2(n1054), .A(n1055), .ZN(n1053) );
  OAI211_X2 U882 ( .C1(n1086), .C2(n1035), .A(n1043), .B(n1087), .ZN(n994) );
  OAI211_X2 U883 ( .C1(in3[2]), .C2(n1034), .A(n431), .B(n428), .ZN(n1087) );
  OAI211_X2 U884 ( .C1(n1069), .C2(n1031), .A(n1038), .B(n1070), .ZN(n1008) );
  OAI211_X2 U885 ( .C1(in4[2]), .C2(n1030), .A(n1040), .B(n491), .ZN(n1070) );
  OAI21_X2 U886 ( .B1(n1071), .B2(n1072), .A(n1073), .ZN(n1040) );
  OAI21_X2 U887 ( .B1(n495), .B2(n493), .A(in4[1]), .ZN(n1073) );
  AOI211_X2 U888 ( .C1(n828), .C2(in4[15]), .A(n829), .B(n830), .ZN(n827) );
  AOI21_X2 U889 ( .B1(n377), .B2(n686), .A(n446), .ZN(n684) );
  OAI21_X2 U890 ( .B1(n1030), .B2(in4[2]), .A(n1031), .ZN(n1029) );
  OAI21_X2 U891 ( .B1(n1034), .B2(in3[2]), .A(n1035), .ZN(n1033) );
  AOI21_X2 U892 ( .B1(n637), .B2(n464), .A(n465), .ZN(n636) );
  AOI21_X2 U893 ( .B1(n642), .B2(n439), .A(n440), .ZN(n641) );
  AOI21_X2 U894 ( .B1(in2[0]), .B2(in4[29]), .A(n549), .ZN(n600) );
  AOI21_X2 U895 ( .B1(n550), .B2(n447), .A(n575), .ZN(n601) );
  AOI21_X2 U896 ( .B1(in1[3]), .B2(in3[25]), .A(n621), .ZN(n663) );
  AOI21_X2 U897 ( .B1(n665), .B2(n443), .A(n444), .ZN(n664) );
  AOI21_X2 U898 ( .B1(in1[1]), .B2(in3[23]), .A(n683), .ZN(n710) );
  AOI21_X2 U899 ( .B1(n712), .B2(n686), .A(n446), .ZN(n711) );
  AOI21_X2 U900 ( .B1(in4[5]), .B2(n1060), .A(n1061), .ZN(n1059) );
  AOI21_X2 U901 ( .B1(in3[21]), .B2(in1[31]), .A(n721), .ZN(n739) );
  OAI21_X2 U902 ( .B1(n740), .B2(n688), .A(n720), .ZN(n738) );
  AOI22_X2 U903 ( .A1(n1054), .A2(in3[5]), .B1(n421), .B2(n425), .ZN(n991) );
  AOI21_X2 U904 ( .B1(in4[21]), .B2(n725), .A(n727), .ZN(n736) );
  OAI21_X2 U905 ( .B1(n737), .B2(n677), .A(n726), .ZN(n735) );
  AOI21_X2 U906 ( .B1(in4[25]), .B2(in2[28]), .A(n613), .ZN(n662) );
  OAI21_X2 U907 ( .B1(n612), .B2(n456), .A(n652), .ZN(n661) );
  OAI211_X2 U908 ( .C1(n615), .C2(n438), .A(n616), .B(n617), .ZN(n556) );
  OAI21_X2 U909 ( .B1(n440), .B2(in1[5]), .A(in3[27]), .ZN(n616) );
  OAI211_X2 U910 ( .C1(n463), .C2(n607), .A(n608), .B(n609), .ZN(n550) );
  OAI21_X2 U911 ( .B1(n465), .B2(in2[30]), .A(in4[27]), .ZN(n608) );
  AOI22_X2 U912 ( .A1(n893), .A2(in4[13]), .B1(n459), .B2(n894), .ZN(n836) );
  AOI22_X2 U913 ( .A1(n398), .A2(in3[13]), .B1(n855), .B2(n887), .ZN(n851) );
  OAI21_X2 U914 ( .B1(n492), .B2(n1039), .A(n1031), .ZN(n1036) );
  OAI21_X2 U915 ( .B1(n1032), .B2(n1044), .A(n1035), .ZN(n1041) );
  AOI211_X2 U916 ( .C1(in2[1]), .C2(n449), .A(n448), .B(n546), .ZN(n545) );
  OAI21_X2 U917 ( .B1(in4[30]), .B2(in2[1]), .A(n550), .ZN(n547) );
  AOI21_X2 U918 ( .B1(n583), .B2(n556), .A(n435), .ZN(n582) );
  OAI21_X2 U919 ( .B1(in3[0]), .B2(n1106), .A(n1089), .ZN(n1105) );
  OAI21_X2 U920 ( .B1(in4[0]), .B2(n1108), .A(n1072), .ZN(n1104) );
  AOI22_X2 U921 ( .A1(in1[27]), .A2(in3[17]), .B1(n412), .B2(n808), .ZN(n760)
         );
  AOI22_X2 U922 ( .A1(in1[31]), .A2(in3[21]), .B1(n380), .B2(n397), .ZN(n689)
         );
  AOI22_X2 U923 ( .A1(n725), .A2(in4[21]), .B1(n470), .B2(n472), .ZN(n679) );
  AOI22_X2 U924 ( .A1(in2[28]), .A2(in4[25]), .B1(n468), .B2(n452), .ZN(n611)
         );
  AOI22_X2 U925 ( .A1(in1[3]), .A2(in3[25]), .B1(n442), .B2(n444), .ZN(n619)
         );
  AOI22_X2 U926 ( .A1(in1[7]), .A2(in3[29]), .B1(n558), .B2(n584), .ZN(n554)
         );
  AOI22_X2 U927 ( .A1(in2[0]), .A2(in4[29]), .B1(n496), .B2(n575), .ZN(n552)
         );
  OAI21_X2 U928 ( .B1(n449), .B2(in2[1]), .A(in4[30]), .ZN(n551) );
  INV_X4 U929 ( .A(reset), .ZN(n1111) );
endmodule

